AM i Wales är oroliga att " framstå som puckon "
Vissa AM , medlemmar i Wales nationalförsamling , är förvirrade över ett förslag att ändra deras titel till MWP ( Member of the Welsh Parliament - Medlem i Wales parlament ) .
Förslaget kommer efter planer på att ändra namnet på nationalförsamlingen till Wales parlament .
AM över hela det politiska spektrumet är oroliga över att bli hånade .
En AM för Labour sa att hans grupp var orolig eftersom " det rimmar med Twp och Pwp " .
För läsare som inte kan walesiska : Twp betyder dum på walesiska och pwp betyder bajs .
En AM för Plaid sa att gruppen i allmänhet var " missnöjd " och har föreslagit andra alternativ .
En konservativ walesare sa att hans grupp är " öppen " för namnändringen , men påpekade att det var ett kort steg från MWP till Mupp .
I det här sammanhanget uttalas W på walesiska likt bokstaven U på engelska i Yorkshire .
Assembly Commission , som för närvarande sammanställer lagstiftning för namnändringen , sa : " Det slutgiltiga beslutet för vad medlemmar i församlingen ska kallas är så klart upp till själva medlemmarna " .
Government of Wales Act 2017 gav den walesiska församlingen rätt att ändra sitt namn .
I juni publicerade kommissionen resultatet av en offentlig konsultation om förslagen , som fann ett starkt stöd för att kalla församlingen för Wales parlament .
Gällande titeln för AM föreslog kommissionen Welsh Parliament Members ( medlemmar i Wales parlament ) eller WMP , men MWP fick störst stöd i en offentlig konsultation .
AM föreslår tydligen andra alternativ , men problem med att nå en konsensus kan orsaka problem för Presiding Officer Elin Jones , som väntas lämna in utkast för lagstiftning om ändringen inom några veckor .
Lagstiftningen för ändringarna inkluderar även andra ändringar för hur församlingen arbetar , inklusive regler för diskvalificering av en AM och utformningen av kommittésystemet .
AM får rösta om vad de ska kallas när de debatterar lagstiftningen .
Makedonien genomför en folkomröstning om ändring av landets namn
På söndag ska väljarna rösta om ifall de ska ändra landets namn till " Republiken Nordmakedonien " .
Folkomröstningen är ett försök att avsluta en dispyt som har pågått i flera årtionden med grannlandet Grekland , som har en provins som heter Makedonien .
Aten har länge insisterat på att grannlandets namn representerar ett anspråk på dess territorium och har upprepade gånger protesterat mot dess försök att bli medlem i EU och NATO .
Makedoniens president Gjorge Ivanov motsätter sig folkomröstningen om namnbytet och har sagt att han kommer att bortse från resultatet .
Men folkomröstningens anhängare , inklusive premiärminister Zoran Zaev , hävdar att namnbytet är priset de måste betala för att gå med i EU och NATO .
Klockorna i St . Martin ' s tystnar när kyrkorna i Harlem stöter på problem
" Äldre personer som jag pratar med säger att det fanns en bar och en kyrka på varje hörn förr " , sa mr Adams .
" Nu finns det varken eller " .
Han sa att det är förståeligt att barerna försvinner .
" Folk umgås på andra sätt nu för tiden " , sa han .
" Barer är inte som områdets vardagsrum längre , dit folk går på regelbunden basis " .
Gällande kyrkorna är han orolig att pengarna från försäljningen av tillgångar inte kommer att räcka så långt som ledarna väntar sig och att " förr eller senare hamnar de på ruta ett igen " .
Han påpekade även att kyrkor kan ersättas av lägenhetsbyggnader med ägarlägenheter fyllda av personer som inte hjälper kvarvarande kyrkor .
" Den absoluta majoriteten av personer som köper lägenheter i byggnaderna kommer att vara vit " , sa han . " Detta kommer så småningom att leda till att alla kyrkorna stängs , eftersom de som flyttar in i lägenheterna förmodligen inte kommer att bli medlemmar i kyrkorna " .
Båda kyrkorna byggdes av vita församlingar innan Harlem blev en svart metropol - Metropolitan Community 1870 , St . Martin ' s ett årtionde senare .
Den ursprungliga vita metodistförsamlingen flyttade ut på 1930 @-@ talet .
En svart församling som hade en kyrka i närheten tog över byggnaden .
St . Martin ' s togs över av en svart församling som leddes av pastor John Howard Johnson , som ledde en bojkott av butiker på 125th Street , en shoppinggata i Harlem , som vägrade anställa eller befordra svarta personer .
Byggnaden skadades allvarligt i en brand 1939 , men när pastor Johnsons församling planerade renoveringen byggde de även klockspelet .
Pastor David Johnson , fader Johnsons son och efterträdare på St . Martin ' s , kallade stolt musikspelet för " de fattigas klockor " .
Experten som spelade klockspelet i juli hade ett annat namn för det : " En kulturell skatt " och " ett oersättligt historiskt instrument " .
Experten , Tiffany Ng från University of Michigan , påpekade även att det var världens första klockspel som spelades av en svart musiker - Dionisio A. Lind , som gick vidare till det större klockspelet i Riverside Church för 18 år sedan .
Enligt mr Merriweather ersatte inte St . Martin ' s honom .
De senaste månadernas händelser på St . Martin ' s är en komplicerad historia med arkitekter och entreprenörer - vissa som anlitats av kyrkans lekmannaskap , andra av det episkopala stiftet .
Kyrkostämman - församlingens styrande organ som består av lekmän - skrev till stiftet i juli och uttryckte en oro för att stiftet skulle " försöka överföra kostnaden " till kyrkostämman , trots att kyrkostämman inte hade varit inblandad när stiftet anlitade arkitekter och entreprenörer .
Vissa församlingsmedlemmar klagade på en brist på transparens från stiftet .
Haj skadar 13 @-@ åring som dyker efter hummer i Kalifornien
I lördags attackerade och skadade en haj en 13 @-@ årig pojke som dök efter hummer i Kalifornien på hummersäsongens första dag , enligt tjänstemän .
Attacken ägde rum strax innan klockan sju på morgonen , nära Beacon ' s Beach i Encinitas .
Chad Hammel sa till KSWB @-@ TV i San Diego att han hade dykt med sina vänner i en halvtimme på lördagsmorgonen när han hörde pojken ropa på hjälp och paddlade dit med en grupp andra för att dra upp honom ur vattnet .
Enligt Hammel trodde han först att pojken bara var glad över att ha hittat en hummer , men sedan insåg han att pojken skrek : " Jag har blivit biten ! "
" Jag har blivit biten ! "
När Hammel kom fram till pojken märkte han att hela nyckelbenen hade slitits upp .
" Jag ropade till alla att ta sig upp ur vattnet . " Det är en haj i vattnet ! " " , berättade Hammel .
Pojken flögs till Rady Children ' s Hospital i San Diego och hans tillstånd anges vara kritiskt .
Det är oklart vilken hajart det var .
Badvaktskaptenen Larry Giles sa till massmedia att en haj hade sett i området några veckor tidigare , men att det hade fastställts att det inte var en farlig hajart .
Giles sa även att offret fick traumaskador på sin övre torso .
Åtkomst till stranden från Ponto Beach i Casablad till Swami ' s i Ecinitas blockerades i 48 timmar av utrednings- och säkerhetsskäl .
Giles nämnde att det finns över 135 hajarter i området , men att de flesta inte anses vara farliga .
Sainsbury ' s ger sig in på Storbritanniens skönhetsmarknad
Sainsbury ' s tar sig an Boots , Superdrug och Debenhams med varuhusliknande skönhetsgångar med skönhetsspecialister .
Som en del av en avsevärd push in i Storbritanniens skönhetsmarknad på £ 2,8 miljarder , som fortsätter växa trots att mode- och hushållsmarknaden faller , kommer de större skönhetsgångarna att testas i 11 butiker landet över och implementeras i fler butiker nästa år om de är framgångsrika .
Investeringen i skönhetsmarknaden är en del av snabbköpens försök att fylla hyllorna som förr togs upp av TV @-@ apparater , mikrovågsugnar och hushållsprodukter .
Sainsbury ' s sa att de tänker fördubbla sitt skönhetsutbud till upp till 3.000 produkter , inklusive märken såsom Revlon , Essie , Tweezerman och Dr . PawPaw för första gången .
Befintliga utbud från L ' Oreal , Maybelline och Burt ' s Bees kommer också att få större utrymme med markerade områden , som i butiker som Boots .
Butikskedjan lanserar även sitt boutique @-@ sminkmärke på nytt så att de flesta av produkterna är veganska - vilket alltfler unga kunder kräver .
Dessutom kommer parfymåterförsäljaren Fragrance Shop att testa stånd i två Sainsbury ' s @-@ butiker - det första ståndet öppnade i Croydon i södra London förra veckan och det andra öppnar i Selly Oak i Birmingham senare i år .
Shopping online och trenden att köpa mindre mängder mat varje dag i lokala butiker innebär att snabbköp måste göra mer för att locka till sig kunder .
Mike Coupe , VD för Sainsbury ' s , har sagt att deras butiker kommer att se ut alltmer som varuhus i ett försök att kämpa emot billiga butiker som Aldi och Lidl med fler tjänster och andra produkter än mat .
Sainsbury ' s har Argos @-@ stånd i hundratals butiker och har även skaffat ett antal Habitat @-@ stånd sedan de köpte båda kedjorna för två år sedan , vilket enligt dem har ökat försäljningen av livsmedel och gjort förvärven lönsammare .
Snabbköpets tidigare försök att ge skönhets- och apoteksavdelningarna ett ansiktslyft misslyckades .
Sainsbury ' s testade ett samarbete med Boots i början av 2000 @-@ talet , men samarbetet avslutades efter en dispyt om hur intäkterna från Boots försäljning i snabbköpen skulle fördelas .
Den nya strategin kommer efter att Sainsbury ' s sålde sin apoteksverksamhet med 281 butiker till Celesio , som äger kedjan Lloyds Pharmacy , för £ 125 miljoner för tre år sedan .
De hävdar att Lloyds skulle spela en roll i planen genom att lägga till ett utökat utbud lyxiga hudvårdsprodukter , inklusive märken som La Roche @-@ Posay och Vichy , i fyra butiker .
Paul Mills @-@ Hicks , Sainsbury ' s kommersiella chef , sa : " Vi har gett våra skönhetsgångar ett nytt utseende och en ny känsla för att förbättra miljön för våra kunder .
Vi har även investerat i särskilt utbildade medarbetare som kan ge kunder råd .
Vårt utbud av märken har utformats för att möta alla behov , och med en tilltalande miljö på smidiga platser är vi nu en lockande skönhetsdestination som utmanar det gamla sättet att shoppa " .
Peter Jones " rasande " efter att Holly Willoughby drar sig ur deal på £ 11 miljoner
Dragons Den @-@ stjärnan Peter Jones är " rasande " över att TV @-@ presentatören Holly Willoughby drar sig ur en deal på £ 11 miljoner med hans livsstilsmärke för att fokusera på sina nya kontrakt med Marks & Spencer och ITV .
Willoughby hinner inte med deras märke Truly , med fritidskläder och tillbehör .
Deras verksamhet har jämförts med Gwyneth Paltrows märke Goop .
This Morning @-@ presentatören , 37 , tillkännagav sitt beslut på Instagram .
Holly Willoughby har gjort Dragons Den @-@ stjärnan Peter Jones rasande genom att dra sig ur deras lukrativa livsstilsmärke i sista minuten - för att fokusera på sina nya avtal med Marks & Spencer och ITV .
Enligt källor blev Jones " rasande " på ett spänt möte på hans affärsimperiums högkvarter i Marlow , Buckinghamshire i tisdags när TV @-@ favoriten medgav att hennes nya avtal - värda upp till £ 1,5 miljon - innebar att hon inte längre hann fokusera på deras märke Truly , med fritidskläder och tillbehör .
Verksamheten har jämförts med Gwyneth Paltrows märke Goop och väntades fördubbla Willoughbys uppskattade förmögenhet på £ 11 miljoner .
När Willoughby , 37 , tillkännagav att hon lämnar Truly på Instagram flög Jones till ett av sina semesterhem .
En källa sa : " Truly var helt klart Hollys främsta prioritet .
Det skulle vara hennes långsiktiga framtid för de kommande årtiondena .
Hennes beslut att dra sig ur chockade alla som var inblandade .
Ingen kunde tro att det hände i tisdags , så nära lanseringen .
Det finns ett lager fullt av varor som är redo att säljas på högkvarteret i Marlow " .
Experter anser att This Morning @-@ presentatörens beslut att dra sig ur kan kosta företaget flera miljoner på grund av avsevärda investeringar i allt från kuddar och ljus till kläder samt risken för vidare förseningar av lanseringen .
Och det kan innebära slutet för en lång vänskap .
Trebarnsmamman Willoughby och hennes man Dan Baldwin har varit nära vänner med Jones och hans fru Tara Capp i tio år .
Willoughby startade Truly med Capp 2016 och Jones , 52 , tog rollen som ordförande i mars .
Paren semestrar tillsammans och Jones äger 40 % av Baldwins TV @-@ produktionsbolag .
Willoughby ska bli märkesambassadör för M & S och kommer att ersätta Ant McPartlin som värd för " I ' m a Celebrity " på ITV .
En källa nära Jones sa i går kväll : " Vi kommenterar inte hans affärsverksamhet " .
Tufft snack " och så blev vi kära "
Han skämtade om att massmedia skulle kritisera honom för en kommentar som vissa skulle anse vara " ovärdig en president " och för att han var så positiv om Nordkoreas ledare .
Varför har president Trump gett upp så mycket ?
Trump sa i en " nyhetsankarröst " :
" Jag har inte gett upp något " .
Han sa att Kim vill ha ett andra möte efter att Trump hyllade deras första möte i Singapore i juni som ett stort steg för Nordkoreas kärnvapennedrustning .
Men förhandlingarna om kärnvapennedrustningen har kört fast .
Mer än tre månader efter mötet i Singapore i juni sa Nordkoreas toppdiplomat Ri Yong Ho till ledarna på FN:s generalförsamling i lördags att Nordkorea inte ser en " motsvarande respons " från USA efter Nordkoreas första nedrustningssteg .
Han noterade att USA i stället fortsätter sanktioner som är avsedda att bibehålla trycket .
Trump var mycket mer optimistisk i sitt tal till sina anhängare .
" Det går jättebra med Nordkorea " , sa han .
" Vi var på väg att kriga med Nordkorea .
Miljontals människor skulle ha dött .
Nu har vi en suverän relation " .
Han sa att hans försök att förbättra relationen till Kim har haft positiva resultat - ett slut på rakettester , befriade gisslan och återlämnade kvarlevor av amerikanska soldater .
Och han försvarade sitt annorlunda sätt att prata om relationen med Kim .
" Det är så lätt att bete sig som en president , men i stället för att ha 10.000 personer som försöker ta sig in i den här fullpackade arenan skulle vi ha runt 200 personer här " , sa Trump och pekade på publiken framför honom .
Tsunami och jordbävning ödelägger ö i Indonesien , hundratals dör
Efter jordbävningen på Lombok , till exempel , blev utländska icke @-@ statliga organisationer tillsagda att de inte behövdes .
Trots att över 10 procent av Lomboks befolkning hade förlorat sina hem utlystes det inte ett undantagstillstånd , vilket krävs för internationellt bistånd .
" I många fall har de tyvärr varit väldigt tydliga med att de inte ber om internationell hjälp , vilket komplicerar det hela " , sa ms Sumbung .
Rädda barnen samlar ett team som ska åka till Palu , men det är ännu oklart om utländsk personal kan arbeta där .
Mr Sutopo , naturkatastrofbyråns talesman , sa att indonesiska tjänstemän utvärderade situationen i Palu för att avgöra om internationella organisationer ska tillåtas delta i biståndsarbetet .
Med tanke på Indonesiens ständiga jordbävningar är landet fortfarande bedrövligt oförberedda på naturens vrede .
Det har byggts tsunamiskydd i Aceh , men de är sällsynta på andra kustlinjer .
Avsaknaden av en tsunamivarningssiren i Palu , trots att en varning hade utfärdats , bidrog förmodligen till förlusten av liv .
Även under perfekta förhållanden är det en utmaning att resa mellan Indonesiens många öar .
Naturkatastrofer komplicerar logistiken ytterligare .
Ett sjukhusfartyg som har legat förankrat i Lombok för att behandla jordbävningsoffer är på väg till Palu , men det tar minst tre dagar för det att nå den nya katastrofen .
President Joko Widodo fokuserade på löften om att förbättra Indonesiens slitna infrastruktur i sin valkampanj och har spenderat stora summor på vägar och tågräls .
Men bristfällig finansiering har plågat mr Jokos administration inför nästa års val .
Mr Joko pressas även av kvardröjande sekteristiska spänningar i Indonesien , där den muslimska majoriteten har antagit en mer konservativ form av tron .
Över 1.000 personer dödades och tiotusentals förlorade sina hem när kristna och muslimska gäng stred på gatorna med machetes , pilbågar och andra primitiva vapen .
Titta på : Liverpools Daniel Sturridge kvitterade i sista minuten mot Chelsea
Daniel Sturridge räddade Liverpool från en Premier League @-@ förlust mot Chelsea med ett mål i 89:e minuten i Stamford Bridge i London i lördags .
Sturridge fick en pass från Xherdan Shaqiri runt 30 meter från Chelseas mål när hans lag låg efter med 1 @-@ 0 .
Han överförde bollen till vänster och scoopade en spark mot den bortre stolpen .
Försöket flög högt över målområdet mot det övre högra hörnet av nätet .
Bollen föll slutligen över Kepa Arrizabalagas hopp och hamnade i nätet .
" Jag försökte bara hamna i en position för att komma åt bollen och spelare som Shaq spelar alltid framåt så mycket som möjligt , så jag försökte bara ge mig själv så mycket tid som möjligt " , sa Sturridge till LiverpoolFC.com.
" Jag såg Kante närma sig och tänkte inte så mycket på det utan sparkade bara " .
Chelsea ledde med 1 @-@ 0 efter första halvleken efter ett mål i 25:e minuten från belgiska stjärnan Eden Hazard .
Den blå strikern hälade en pass tillbaka till Mateo Kovacic , spinnade av nära mittfältet och sprintade till Liverpools sida .
Kovacic gjorde en snabb give @-@ and @-@ go vid mittfältet .
Sedan fick han en suverän spark som förde in Hazard i målområdet .
Hazard sprang ifrån försvaret och fick bollen i nätet vid den bortre stolpen med en vänsterfotad spark förbi Liverpools Alisson Becker .
Liverpool kämpar mot Napoli i gruppstadiet av Champions League på Stadio San Paolo i Neapel , Italien klockan 15 : 00 på onsdag .
Chelsea ställs emot VIdeoton i Uefa Europa League i London klockan 15 : 00 på torsdag .
Dödssiffra för tsunami i Indonesien stiger till 832
Dödssiffran för jordbävningen och tsunamin i Indonesien har stigit till 832 , enligt landets katastrofbyrå tidigt i söndags .
Många människor rapporterades ha fastnat i spillrorna av byggnader som rasat i jordbävningen på 7,5 som slog till i fredags och utlöste vågor på upp till sex meter , sa byråns talesman Sutopo Purwo Nugroho på en nyhetskonferens .
Staden Palu , med över 380.000 invånare , var full av bråte från byggnader som rasat .
Polisen griper man , 32 , misstänkt för mord efter att kvinna huggs ihjäl
En mordutredning har startats efter att en kvinnas lik hittades i Birkenhead , Merseyside i morse .
44 @-@ åringen hittades klockan 7 : 55 med knivsår på Grayson Mews på John Street , och en 32 @-@ årig man greps misstänkt för mord .
Polisen har bett personer i området som såg eller hörde något att träda fram .
Kriminalinspektör Brian O ' Hagan sa : " Vi är i ett tidigt stadium av utredningen , men jag ber alla som var i närheten av John Street i Birkenhead och såg eller hörde något misstänkt att kontakta oss .
Jag ber även alla , särskilt taxiförare , som kan ha filmat något med en bilkamera att kontakta oss eftersom de kan ha information som är avgörande för vår utredning " .
En talesman för polisen har bekräftat att kvinnan som hittades bor i Birkenhead och att kroppen hittades inuti en fastighet .
Under eftermiddagen har vänner som tror att de känner kvinnan anlänt till platsen för att fråga var hon hittades i morse .
Utredningen pågår och polisen underrättar offrets närmaste anhörige .
En taxiförare som bor i Grayson Mews har precis försökt komma in i sin lägenhet , men polisen sa att ingen får komma in i eller gå ut ur byggnaden .
Han blev mållös när han fick reda på vad som hade hänt .
De boende i byggnaden har underrättats om att det tar flera timmar innan de får komma in igen .
En polisassistent sa till en man att hela området behandlas som en brottsplats .
En gråtande kvinna dök upp på platsen .
Hon säger " det är så hemskt " om och om igen .
Klockan 14 : 00 stod det två polisbilar innanför avspärrningen och en annan precis utanför .
Ett antal polisassistenter stod innanför avspärrningen med översikt över lägenhetsbyggnaden .
Personer med information ombes skicka ett DM till @ MerPolCC , ringa 101 eller kontakta Crimestoppers anonymt på 0800 555 111 och ange logg 247 från 30 september .
Parlamentets staty av Cromwell senaste offer för gräl om omskrivning av historien
En bannlysning vore poetisk rättvisa för hans talibanliknande förstörelse av så många av Englands kulturella och religiösa artefakter som utfördes av hans fanatiska puritanska följare .
Men Cromwell Society kallade mr Cricks förslag för " dårskap " och " försök att skriva om historien " .
John Goldsmith , ordförande för Cromwell Society , sa : " Det var oundvikligt att statyn av Oliver Cromwell utanför Westminsterpalatset skulle dras in i den pågående debatten om att ta bort statyer " .
Ikonoklasmen under de engelska inbördeskrigen varken beordrades eller utfördes av Cromwell .
Fel Cromwell kanske skulle offras för det hans förfader Thomas gjorde 100 år tidigare .
Sir William Hamo Thorneycrofts magnifika representation av Cromwell visar 1800 @-@ talets åsikt om och är en del av historiografin för en man som många anser fortfarande bör hyllas .
Mr Goldsmith sa till The Sunday Telegraph : " Många , kanske fler på slutet av 1800 @-@ talet än nu , anser att Cromwell försvarade parlamentet mot tryck utifrån , i hans fall från monarkin .
Om detta är en korrekt representation är föremål för en pågående historisk debatt .
Men konflikten under mitten av 1600 @-@ talet har utan tvekan påverkat vår nations utveckling , och Cromwell är en välkänd person som representerar ena sidan av saken .
Hans bedrifter som lordprotektor förtjänar också att hyllas och firas .
Mördargris dödar bonde
En bonde attackerades och dödades av en gris på en marknad i sydvästra Kina , enligt lokala mediarapporter .
Mannen , som endast identifieras med sitt efternamn Yuan , hittades död med en brusten artär och täckt i blod i en stia på marknaden i Liupanshui i provinsen Guizhou , rapporterade South China Morning Post i söndags .
En grisuppfödare gör sig redo att injicera vaccin i grisar i en svinstia den 30 maj 2005 i Xining i provinsen Qinghai , Kina .
Han rapporteras ha färdats med sin kusin från grannprovinsen Yunnan i onsdags för att sälja 15 grisar på marknaden .
Morgonen därpå hittade kusinen honom död och upptäckte att dörren till en svinstia i närheten var öppen .
Han sa att det fanns en stor grishane i svinstian med blod på munnen .
En rättsteknisk undersökning bekräftade att den 250 kilo tunga grisen hade dödat bonden , enligt rapporten .
" Min kusins ben var blodiga och förvridna " , sa kusinen som identifieras med efternamnet Wu till Guiyang Evening News .
En övervakningskamera filmade Yuan när han kom till marknaden för att mata sina grisar klockan 4 : 40 i torsdags .
Hans kropp hittades en timme senare .
Grisen som dödade bonden tillhörde inte Yuan eller hans kusin .
En marknadsmanager sa till Evening News att grisen hade låsts in för att undvika fler attacker medan polisen samlade in bevis på platsen .
Yuans familj och de ansvariga för marknaden rapporteras förhandla om kompensation för hans död .
Det är sällsynt att grisar attackerar människor , men det har hänt förut .
2016 attackerade en gris en kvinna och hennes man på deras gård i Massachusetts och gav mannen allvarliga skador .
Tio år tidigare tryckte en gris på 300 kilo fast en bonde i Wales mot en traktor tills hans fru skrämde bort den .
När en bonde i Oregon blev uppäten av sina grisar 2012 sa en bonde i Manitoba till CBC News att grisar normalt sett inte är aggressiva , men att smaken av blod kan fungera som en " katalysator " .
" De är bara lekfulla .
De nafsar och är väldigt nyfikna . De vill inte skada någon .
Man måste bara visa dem respekt " , sa han .
Resterna av orkanen Rosa för vidsträckt kraftigt regn till sydvästra USA
Som förutsett blir orkanen Rosa svagare när den färdas över svalare vatten vid Mexikos norra kust .
Men Rosa kommer att föra med sig översvämmande regn till norra Mexiko och sydvästra USA de kommande dagarna .
Rosa hade en vindstyrka på upp till 135 km / tim , kategori 1 , klockan fem EST i söndags och befann sig 620 km sydväst om Punta Eugenia , Mexiko .
Rosa väntas färdas norrut på söndag .
Under tiden börjar en tråg bildas över Stilla havet och färdas österut mot USA:s västra kust . När Rosa närmar sig halvön Baja California som en tropisk storm på måndag kommer den att tvinga djup tropisk fukt norrut in i sydvästra USA .
Rosa kommer att föra med sig upp till 25 cm regn i vissa delar av Mexiko på måndag .
Sedan kommer tropisk fukt som interagerar med den närmande trågen att skapa vidsträckt kraftigt regn i sydvästra USA de kommande dagarna .
Lokalt kommer 2,5 @-@ 10 cm regn att orsaka farlig översvämning , lerflöden och möjligen jordskred i öknen .
Djup tropisk fukt kommer att leda till 5 @-@ 7,5 cm regn per timme på vissa platser , särskilt i delar av södra Nevada och Arizona .
Upp till 5 @-@ 10 cm regn väntas på vissa platser i sydvästra USA , särskilt i stora delar av Arizona .
Plötsliga översvämningar är möjliga med snabbt försämrade förhållanden på grund av det utspridda tropiska regnet .
Det rekommenderas absolut inte att någon ger sig ut i öknen till fots när tropiskt regn väntas .
Kraftigt regn kan göra kanjoner till forsande floder och åskstormar leder till starka lokala vindar som blåser runt sand .
Den närmande trågen för med sig visst lokalt kraftigt regn till delar av södra Kaliforniens kustlinje .
Det är möjligt med sammanlagt över en cm regn , vilket kan leda till lerflöden och hala vägar .
Det vore det första regnet i området under regnperioden .
Vissa skingrade tropiska regnskurar kommer att närma sig Arizona sent på söndag och tidigt på måndag , innan regnet blir mer vidsträckt senare på måndagen och tisdagen .
Kraftigt regn kommer att spridas till Four Corner på tisdag och fortsätta under onsdagen .
Oktober kan innebära intensiva temperaturförändringar i hela USA , när Arktis kyls ned men tropikerna förblir varma .
Ibland leder detta till dramatiska temperaturförändringar på korta avstånd .
Det finns ett bra exempel på dramatiska temperaturskillnader i centrala USA på söndag .
Det är nästan tio graders skillnad mellan Kansas City i Missouri och Omaha i Nebraska , och mellan St . Louis och Des Moines i Iowa .
Under de kommande dagarna kommer den kvarvarande sommarvärmen att försöka spridas igen .
Stora delar av centrala och östra USA väntas få en varm start på Oktober med runt 30 grader från Great Plains till delar av nordöstra USA .
New York kan få 27 grader på tisdag , vilket vore runt fem grader över genomsnittet .
Vår långsiktiga klimatprognos tyder på stor chans för varmare temperaturer än genomsnittet i östra USA under första halvan av oktober .
Över 20 miljoner tittade på Brett Kavanaughs förhör
Över 20 miljoner tittade på torsdagens gripande vittnesmål från Brett Kavanaugh , som nominerats till högsta domstolen , och Christine Blasey Ford , som anklagade honom för sexuellt överfall som ska ha ägt rum på 1980 @-@ talet , på sex TV @-@ nätverk .
Under tiden fortsatte det politiska dödläget och den normala sändningen avbröts för fredagens sista minuten @-@ twist - Arizonas senator Jeff Flakes avtal med FBI där de fick en vecka på sig att utreda anklagelsen .
Ford sa till Senate Judiciary Committee att hon är helt säker på att Kavanaugh tafsade på henne när han var full och försökte ta av hennes kläderna på en high school @-@ fest .
Kavanaugh gav ett passionerat vittnesmål och sa att han är helt säker på att det inte hände .
Det är troligt att antalet tittare i fredags var högre än de 20,4 miljoner som angetts av Nielsen .
De räknade genomsnittligt antal tittare på CBS , ABC , NBC , CNN ; Fox News Channel och MSNBC .
Antalet tittare var inte omedelbart tillgängligt för andra TV @-@ nätverk som visade förhöret , inklusive PBS , C @-@ SPAN och Fox Business Network .
Och Nielsen har ofta problem att räkna personer som tittar från kontor .
Jämförelsevis är det lika många tittare som för en footballmatch i slutspelet eller Oscarsgalan .
Fox News Channel , vars presentatörer har visat ett starkt stöd för Kavanaughs nominering , hade flest tittare med ett genomsnitt på 5,69 miljoner under det dagslånga förhöret , enligt Nielsen .
ABC hade näst flest med 3,26 miljoner tittare .
CBS hade 3,1 miljon , NBC hade 2,94 miljoner , MSNBC hade 2,89 miljoner och CNN hade 2,52 miljoner , enligt Nielsen .
Intresset var fortsatt högt efter förhöret .
Flake var i fokus under fredagens drama .
Efter att republikanens kontor utfärdade ett uttalande om att han skulle rösta för Kavanaugh filmade CNN och CBS demonstranter som skrek på honom när han försökte ta en hiss till ett förhör med Judiciary Committee på fredagsmorgonen .
Han tittade ned på golvet i flera minuter medan demonstranterna skrek på honom , vilket visades i direktsändning av CNN .
" Jag står ju rakt framför dig " , sa en kvinna .
Tror du att han berättar sanningen för landet ? "
De sa även : " Du har makt när så många kvinnor är maktlösa " .
Flake sa att hans kontor hade utfärdat ett uttalande och innan hissdörrarna stängdes sa han att han skulle ha mer att säga efter förhöret med kommittén .
TV @-@ nätverken sände live flera timmar senare när Judiciary Committee röstade om ifall de skulle föra vidare Kavanaughs nominering till en omröstning med hela senaten .
Men Flake sa att han endast tänkte göra det om FBI skulle utreda anklagelserna mot den nominerade under den kommande veckan , vilket minoritetsdemokraterna har yrkat på .
Flake blev delvis övertygad av sin vän , den demokratiska senatorn Chris Coons .
Efter att ha pratat med Coons och flera senatorer efteråt fattade Flake sitt beslut .
Flakes beslut hade stor påverkan , eftersom det var tydligt att republikanerna inte skulle ha tillräckligt med röster för att godkänna Kavanaugh utan utredningen .
President Trump har startat en FBI @-@ utredning om anklagelserna mot Kavanaugh .
Brittiska premiärministern May anklagar kritiker för " politiska lekar " kring Brexit
Premiärminister Theresa May har anklagat kritiker av hennes planer om att lämna Europeiska unionen för " politiska lekar " om Storbritanniens framtid och att underminera nationens intresse i en intervju med tidningen Sunday Times .
Storbritanniens premiärminister Theresa May anländer till den konservativa partikonferensen i Birmingham , Storbritannien 29 september 2018 .
I en annan intervju bredvid hennes på tidningens framsida fortsatte hennes före detta utrikesminister Boris Johnson sin attack mot hennes så kallade Chequers @-@ plan för Brexit och sa att förslaget om att Storbritannien och EU ska samla in varandras tullavgifter var " fullständigt orimligt " .
Skjutningen av Wayde Sims : Polisen griper misstänkte Dyteon Simpson för LSU @-@ spelarens död
Polisen har gripit en misstänkt för dödsskjutningen av Wayde Sims , en 20 @-@ årig basketspelare på LSU .
Dyteon Simpson , 20 , har gripits och satts i häktet för mord , sa polisen i Baton Rouge .
Myndigheterna släppte en video av konfrontationen mellan Sims och Simpson och polisen sa att Sims tappade sina glasögon i striden .
Polisen hittade glasögonen på platsen och fann Simpsons DNA på dem , enligt CBS dotterbolag WAFB .
Efter förhör med Simpson sa polisen att han erkände att han sköt ihjäl Wayde .
Hans borgen fastställdes till 350.000 dollar , enligt Advocate .
Rättsläkaren i East Baton Rouge Parish släppte en preliminär rapport i fredags , enligt vilken dödsorsaken var ett skottsår i huvudet och in i nacken .
Polisen tackar Louisiana State Polices rymlingsinsatsstyrka , polisens statliga rättslabb , Southern Universitys polis och invånare i området för hjälp med utredningen som ledde till gripandet .
LSU:s atletiska direktör Joe Alleva tackade den lokala polisen för deras " flit och strävan efter rättvisa " .
Sims var 20 år .
Den 1,98 meter långa forwarden växte upp i Baton Rouge , där hans pappa Wayne också spelade basket för LSU .
Han hade ett genomsnitt på 5,6 poäng och 2,6 rebounds per match förra säsongen .
I fredags morse sa LSU:s baskettränare Will Wade att laget var " förkrossat " och " chockat " av Waydes död .
" Man är orolig för sådant här hela tiden " , sa Wade .
Vulkan spyr aska över Mexico City
Aska från vulkanen Popocatépetl har nått den södra delen av Mexikos huvudstad .
National Center for Disaster Prevention varnade i lördags mexikaner att hålla sig borta från vulkanen efter att aktivitet hade upptäckts i kratern och de registrerade 183 utsläpp av gas och aska under loppet av 24 timmar .
Centret upptäckte flera muller och skalv .
Bilder på sociala medier visade tunna lager av aska på vindrutor i områden av Mexico City , som Xochimilco .
Geofysiker har noterat ökad aktivitet i vulkanen som står 72 km sydost om huvudstaden sedan en jordbävning på 7,1 drabbade centrala Mexiko i september 2017 .
Vulkanen som kallas Don Goyo har varit aktiv sedan 1994 .
Polis drabbar samman med katalanska separatister inför årsdagen för självständighetsomröstningen
Sex personer greps i Barcelona i lördags efter att självständighetsdemonstranter drabbade samman med kravallpolis samtidigt som tusentals personer deltog i rivaliserande demonstrationer för att markera den första årsdagen för Kataloniens polariserande omröstning om secession .
En grupp maskerade separatister som hölls tillbaka av kravallpolis kastade ägg och färgpulver på dem , vilket ledde till mörka dammoln på gator som i vanliga fall är fulla av turister .
Slagsmål bröt även ut senare under dagen och poliser använde sina batonger för att stoppa dem .
Under flera timmar ropade självständighetsgrupperna " aldrig glömma , aldrig förlåta " medan unionisterna ropade " länge leve Spanien " .
14 personer behandlades för mindre skador som orsakats av protesterna , enligt lokal press .
Stämningen är fortfarande spänd i regionen som längtar efter självständighet ett år efter folkomröstningen den första oktober som ansågs vara illegal av Madrid men hyllades av katalanska separatister .
En överväldigande majoritet röstade för självständighet , men deltagandet var lågt då de flesta som var emot secessionen bojkottade omröstningen .
Enligt katalanska myndigheter skadades nästan 1.000 personer i våldsamma sammandrabbningar i fjol när polisen försökte stoppa omröstningen vid valstationer i regionen .
Självständighetsgrupper campade under natten på fredagen för att förhindra en demonstration till stöd för den nationella polisen .
Demonstrationen ägde rum ändå , men tvingades ta en annan rutt .
Elektrikern Narcis Termes , 68 , deltog i separatisternas protest med sin fru och sa att han inte längre tror att Katalonien kommer att bli självständigt .
" I fjol upplevde vi en av våra bästa stunder .
Jag såg mina föräldrar gråta av glädje över att kunna rösta , men nu har vi kört fast " , sa han .
Trots en avgörande men marginal vinst i regionala val i december har katalanska partier som är för självständigheten haft svårt att hålla drivkraften uppe i år , då många av deras mest välkända ledare lever i självpålagd exil eller sitter i häkte i väntan på rättegång om deras roll i organiseringen av folkomröstningen och den efterföljande självständighetsförklaringen .
Joan Puig , en 42 @-@ årig mekaniker som spelade in protesten till stöd för polisen på sin mobil , sa att konflikten hade fyrats på av politiker på båda sidor .
" Det blir alltmer spänt " , sa han .
I lördags tillkännagav Oriol Junqueras , en av nio katalanska ledare som har suttit i häkte sedan i slutet av förra året , att han tänker kandidera i valet till Europaparlamentet nästa år .
" Att kandidera till Europaparlamentet är det bästa sättet att fördöma återgången av demokratiska värderingar och det underkuvande vi har upplevt från den spanska regeringen " , sa han .
Londonderry : Män gripna efter att bil kör in i hus
Tre män - 33 , 34 och 39 - har gripits efter att en bil kördes in i ett hus i Londonderry upprepade gånger .
Incidenten ägde rum i Ballynagard Crescent , runt klockan 19 : 30 BST i torsdags .
Kriminalinspektör Bob Blemmings sa att grindarna och själva byggnaden skadades .
En armborst kan även ha avfyrats mot bilen .
Menga ger Livingston 1 @-@ 0 mot Rangers
Dolly Mengas första mål för Livingston säkrade vinsten
Livingston chockade Rangers och dömde Steven Gerrard till sin andra förlust på 18 matcher som manager för Ibrox @-@ klubben .
Dolly Mengas strike visade sig vara skillnaden när Gary Holts sida blev delad tvåa med Hibernian .
Gerrards sida har fortfarande inte fått en bortavinst i Premiership den här säsongen och möter Hearts , med åtta poäng mer , nästa söndag .
Innan dess välkomnar Rangers Rapid Vienna i Europa League på torsdag .
Livingston förlänger sin vinststräcka till sex matcher - huvudtränaren Holt har fortfarande inte upplevt en förlust sedan han ersatte Kenny Miler förra månaden .
Livingston missar chanser mot tvära besökare
Holts lag borde ha tagit ledningen långt innan de gjorde mål ; deras rättframhet gav Rangers alla möjliga problem .
Scott Robinson bröt sig igenom men släpade sin prestation tvärs över målet , och sedan kunde Alan Lithgow bara skjuta brett efter att ha glidit in för att mäta Craig Halketts nickning tvärs över målet .
Hemmalaget nöjde sig med att låta Rangers spela framför dem , då de visste att de kunde attackera i bestämda spel .
Och det var så det avgörande målet gjordes .
Rangers gav upp en frispark och Livingston utnyttjade en öppning . Declan Gallagher och Robinson samarbetade för att ge Menga en chans , som gjorde mål från mitten av målområdet .
I det läget hade Rangers dominerat bollen , men hemmalagets försvar var ogenomträngligt och målvakten Liam Kelly lämnades i stort sett i fred .
Samma mönster fortsatte i andra halvleken , men Alfredo Morelos tvingade fram en räddning från Kelly .
Scott Pittman nekades av Rangers målvakt Allan McGregors fötter och Lithgow sköt brett från en annan av Livingstons bestämda spel .
Korsningar kom ständigt in i Livingstons målområde och hanterades utan problem . Två straffkrav - efter Halketts utmaning av utbytaren Glenn Middleton och en för hands - avfärdades .
" Fenomenal " från Livingston - analys
BBC Scotlands Alasdair Lamont på Tony Macaroni Arena
Fenomenal uppvisning och resultat för Livingston .
Varenda en var enastående och fortsätter överskrida förväntningarna på vägen uppåt .
Deras spelstil och personal har knappt förändrats sedan de återvände till övre nivån , men Holt förtjänar äran för att ha galvaniserat laget sedan sin ankomst .
Han hade så många hjältar .
Kapten Halkett var enastående och ledde ett skickligt organiserat försvar , och Menga höll Connor Goldson och Joe Worrall på helspänn rakt igenom .
Men Rangers saknade inspiration .
De har haft sina stunder under Gerrard , men de levde inte upp till standarden .
Deras sista boll höll inte måttet - de öppnade bara hemmasidan en gång - och det är något av en väckarklocka för Rangers , som ligger i mitten .
Erdogan får ett blandat välkomnande i Köln
Lördagen bjöd på leenden och blå himmel ( 29 september ) när Turkiets och Tysklands ledare åt frukost tillsammans i Berlin .
Det är den sista dagen av president Erdogans kontroversiella besök i Tyskland - som ska reparera relationen mellan de NATO @-@ allierade .
De har blivit osams över mänskliga rättigheter , tryckfrihet och Turkiets inträde i EU .
Erdogan åkte sedan till Köln för att öppna en enorm ny moské .
Staden har världens största turkiska befolkning utanför Turkiet .
Polisen hävdade att de hindrade 25.000 åskådare från att samlas utanför moskén av säkerhetsskäl , men många anhängare samlades i närheten för att se sin president .
Hundratals anti @-@ Erdogan @-@ demonstranter - många av dem kurdiska - gjorde även sina röster hörda och fördömde både Erdogans policyer och den tyska regeringens beslut att välkomna honom till Tyskland .
De duellerande protesterna visar de splittrade åsikterna om en besökare som anses vara en hjälte av vissa tyska turkar och fördöms som en envåldshärskare av andra .
Vägolycka i Deptford : Cyklist dör i krock med bil
En cyklist har dött i en krock med en bil i London .
Krocken ägde rum nära korsningen av Bestwood Street och Evelyn Street , en vältrafikerad väg i Deptford i sydöstra London , runt klockan 10 : 15 BST .
Bilföraren stannade bilen och sjukvårdare kallades dit , men mannen dog på platsen .
Krocken äger rum några månader efter att en annan cyklist dog i en smitningsolycka på Childers Street , runt 1,5 km från krocken i lördags .
Metropolitan Police sa att de försöker identifiera mannen och underrätta hans närmaste anhöriga .
Vägar har spärrats av och bussar har omdirigerats och bilförare ombeds undvika området .
Long Lartin @-@ fängelset : Sex vakter skadade i tumult
Sex fängelsevakter har skadats i oroligheter på ett högsäkerhetsfängelse för män , enligt Prison Office .
Oroligheterna bröt ut på HMP Long Lartin i Worcestershire runt klockan 9 : 30 BST i söndags och pågår fortfarande .
Specialiserade " tornadovakter " har kallats dit för att hantera oroligheterna , som involverar åtta fångar på en flygel .
Vakterna behandlades på plats för smärre skador i ansiktet .
En talesperson för Prison Service sa : " Särskilt utbildad fängelsepersonal har skickats dit för att hantera den pågående incidenten på HMP Long Lartin .
Sex personalmedlemmar har behandlats för skador .
Vi tolererar inte våld i våra fängelser och är tydliga med att de som ligger bakom detta kommer att hänföras till polisen och kan få utökade fängelsestraff " .
HMP Long Lartin rymmer över 500 fångar , inklusive några av landets farligaste förbrytare .
I juni rapporterades det att fängelsets direktör behandlades på sjukhus efter att ha blivit attackerad av en fånge .
Och i oktober i fjol kallades kravallpolis till fängelset för att hantera allvarliga oroligheter där personal attackerades med biljardbollar .
Orkanen Rosa hotar Phoenix , Las Vegas , Salt Lake City med översvämning ( områden med torka kan dra nytta )
Det är sällsynt att tropiska lågtryck når Arizona , men det är precis vad som troligen kommer att hända i början av nästa vecka när orkanen Rosas kvarvarande energi drar fram över öknen i sydvästra USA , med risk för plötslig översvämning .
National Weather Service har redan utfärdat varningar för plötsliga översvämningar för måndag och tisdag i västra Arizona och in i södra och östra Nevada , sydöstra Kalifornien och Utah , inklusive städerna Phoenix , Flagstaff , Las Vegas och Salt Lake City .
Rosa väntas färdas direkt över Phoenix på tisdag , och föra med sig regn sent på måndag .
National Weather Service i Phoenix sa i ett tweet att endast " tio tropiska cykloner har bibehållit status som tropisk storm eller lågtryck inom 320 km från Phoenix sedan 1950 !
Katrina ( 1967 ) var en orkan inom 65 km från Arizonas gräns " .
National Hurricane Centers senaste modeller förutspår 5 @-@ 10 cm regn , med isolerade mängder på upp till 15 cm i Mogollon Rim i Arizona .
Andra delar av öknen i sydvästra USA , inklusive centrala Klippiga bergen och Great Basin , får förmodligen 2,5 @-@ 5 cm regn med risk för upp till 10 cm .
I områden utan risk för plötsliga översvämningar kan Rosas regn vara en välsignelse , eftersom regionen är drabbad av torka .
Översvämningar är väldigt allvarliga , men en del av regnet kommer förmodligen att vara till nytta eftersom sydvästra USA lider av torka .
Enligt U.S. Drought Monitor lider strax över 40 procent av Arizona av åtminstone extrem torka , den näst högsta kategorin , rapporterade weather.com.
Orkanen Rosa kommer först att färdas över halvön Baja California i Mexiko .
Rosa , fortfarande med orkanstyrka i söndags morse med maxvindstyrka på 135 km / tim , befinner sig 620 km söder om Punta Eugenia i Mexiko och färdas norrut i 20 km / tim .
Stormen stöter på svalare vatten i Stilla havet , vilket lugnar ned den .
Den väntas därför nå Mexikos landmassa som en tropisk storm på måndag eftermiddag eller kväll .
Delar av Mexiko kan få kraftigt regn , vilket utgör en avsevärd risk för översvämning .
" Sammanlagt 7,5 @-@ 15 cm regn väntas från Baja California till nordvästra Sonora , med en risk för upp till 25 cm " , rapporterade weather.com.
Rosa kommer sedan att färdas norrut över Mexiko som en tropisk storm och nå Arizonas gräns tidigt tisdag morgon som ett tropiskt lågtryck , som sedan kommer att färdas genom Arizona och in i södra Utah sent tisdag kväll .
" Den största faran från Rosa och dess kvarvarande energi är väldigt kraftigt regn i Baja California , nordvästra Sonora och öknen i sydvästra USA " , sa National Hurricane Center .
Regnet väntas leda till livshotande plötsliga översvämningar och lerflöden i öknen , samt jordskred i bergig terräng .
Attack i Midsomer Norton : Fyra gripna för mordförsök
Tre pojkar i tonåren och en 20 @-@ årig man har gripits misstänkta för mordförsök efter att en 16 @-@ åring hittades med knivsår i Somerset .
Den tonåriga pojken hittades skadad i området Excelsior Terrace i Midsomer Norton , runt klockan 4 : 00 BST i lördags .
Han togs till sjukhus och läget rapporteras vara " stabilt " .
En 17 @-@ åring , två 18 @-@ åringar och en 20 @-@ årig man greps under natten i området Radstock , sa polisen i Avon och Somerset .
Polisen ber alla som kan ha filmat det som hände med mobilen att träda fram .
Trump säger att Kavanaugh " led , elakheten , ilskan " från demokratiska partiet
" En röst för domare Kavanaugh är en röst för att förkasta det demokratiska partiets hänsynslöshet och skandalösa taktiker " , sa Trump till sina anhängare i Wheeling , West Virginia .
Trump sa att Kavanaugh hade " lidit av elakheten , ilskan " från det demokratiska partiet under hela nomineringsprocessen .
Kavanaugh vittnade inför kongressen i torsdags och förnekade starkt och känslosamt Christine Blasey Fords anklagelse att han förgrep sig sexuellt på henne flera årtionden tidigare då de var tonåringar .
Ford vittnade också inför kongressen om sin anklagelse .
Presidenten sa i lördags att " det amerikanska folket såg det briljanta och kvaliteten och modet " hos Kavanaugh den dagen .
" En röst för att bekräfta domare Kavanaugh är en röst för att bekräfta en av våra tiders skickligaste juridiska sinnen , en jurist med en förstklassig historia av att tjäna allmänheten " , sa han till sina anhängare i publiken i West Virginia .
Presidenten hänvisade indirekt till Kavanaughs nominering när han pratade om vikten av att republikaner röstar i de kommande midterm elections .
" Vi är fem veckor från ett av våra livs viktigaste val .
Jag kandiderar inte , men jag kandiderar " , sa han .
" Det är därför jag åker runt och kämpar för suveräna kandidater " .
Trump hävdade att demokraterna försöker " stå emot och hindra " .
Den första avgörande omröstningen i senaten om Kavanaughs nominering väntas äga rum senast fredag , enligt information till CNN från en assistent till en senior republikansk ledare .
Hundratals döda i jordbävning och tsunami i Indonesien , antalet stiger
Minst 384 personer dog , många sveptes bort när gigantiska vågor kraschade mot stränderna , när en stor jordbävning och tsunami drabbade den indonesiska ön Sulawesi , enligt myndigheterna i lördags .
Hundratals personer hade samlats för en festival på stranden i staden Palu i fredags när upp till sex meter höga vågor kraschade mot stranden i skymningen och svepte ut många till en säker död och förstörde allt i sin väg .
Tsunamin kom efter en jordbävning på 7,5 .
" När tsunamivarningen kom i går stannade folk på stranden i stället för att omedelbart springa därifrån , och de föll offer för tsunamin " , sa Sutopo Purwo Nugroho , talesman för Indonesiens katastrofbyrå BNPB , på ett möte i Jakarta .
" Tsunamin var inte ensam utan släpade med sig bilar , stockar och hus . Den drabbade allt i dess väg " , sa Nugroho . Han sa även att tsunamin hade färdats på öppet hav i upp till 800 km / tim innan den drabbade kustlinjen .
En del klättrade upp i träd för att komma undan tsunamin och överlevde , sa han .
Runt 16.700 personer evakuerades till 24 anläggningar i Palu .
Flygfoton som släppts av katastrofbyrån visar att många byggnader och butiker är förstörda , broar är förvridna och har kollapsat och en moské är omgiven av vatten .
Efterskalv drabbade fortfarande kuststaden i lördags .
Raden av jordbävningar kändes i ett område med en befolkning på 2,4 miljoner .
Indonesiens byrå för utvärdering och tillämpning av teknik BPPT sa i ett uttalande att den mängd energi som frigjordes i den enorma jordbävningen i fredags var 200 gånger så stor som atombomben som släpptes på Hiroshima i andra världskriget .
Staden ligger i änden av en lång , smal bukt , vilket kan ha gjort tsunamin större , enligt byrån .
Nugroho beskrev förödelsen som " omfattande " och sa att tusentals hus , sjukhus , köpcenter och hotell har kollapsat .
Döda offer hittades under bråtet av kollapsade byggnader , sa han , och 540 personer skadades och 29 är saknade .
Nugroho sa att offren och skadorna kan vara ännu värre längs kustlinjen 300 km norr om Palu , ett område som kallas Donggala , som är närmre jordbävningens epicenter .
Kommunikationen från Donggala " var helt förlamad utan någon information " , sa Nugroho .
" Det bor över 300.000 personer där " , sa Röda korset i ett uttalande , och dess personal och volontärer är på väg till de drabbade områdena .
" Det är redan en tragedi , men det kan bli mycket värre " , sa de .
Byrån kritiserades i lördags för att inte ha informerat om att tsunamin hade slagit till mot Palu , men myndigheterna sa att vågorna hade dykt upp inom tiden som varningen utfärdades .
I en amatörvideo som delats på sociala medier hörs en man på övervåningen i en byggnad skrika frenetiska varningar om tsunamin till personer på gatan nedanför .
Inom några minuter kraschar en mur av vatten mot stranden och sveper bort byggnader och bilar .
Reuters kunde inte omedelbart autentisera videon .
Jordbävningen och tsunamin ledde till ett omfattande strömavbrott som avbröt all kommunikation runt Palu , vilket försvårade räddningsarbetet för myndigheterna .
Militären har börjat skicka dit lastflyg med hjälp från Jakarta och andra städer , enligt myndigheterna , men evakuerade personer är fortfarande i stort behov av mat och andra förnödenheter .
Stadens flygplats har öppnats för hjälparbetet och förblir stängd för övrig trafik till oktober .
President Joko Widodo planerade att besöka anläggningar i Palu på söndag .
Antalet döda i tsunami i Indonesien överstiger 800 .
Det är väldigt illa .
Medarbetare från World Vision i Donggala har tagit sig till Palu där de söker skydd under presenningar på gården utanför kontoret , men de såg förödelse längs vägen , enligt mr Doseba .
" De sa att de såg många förstörda hus " , sa han .
Det är väldigt illa .
Biståndsgrupper har påbörjat det bistra biståndsarbetet , men vissa klagade på att utländska biståndsarbetare med omfattande expertis hindrades från att resa till Palu .
Enligt indonesiska föreskrifter får finansiering , förnödenheter och medarbetare från utomlands endast användas om undantagstillstånd utlyses efter en katastrof .
Detta har ännu inte hänt .
" Det är fortfarande en regional katastrof " , sa Aulia Arriani , en talesperson för indonesiska Röda korset .
" När myndigheterna säger att det är en nationell katastrof kan vi släppa in internationellt bistånd , men den statusen har inte utlysts än " .
När den andra kvällen föll i Palu efter fredagens jordbävning och tsunami hoppades släkt och vänner till saknade personer fortfarande på att deras nära och kära skulle visa sig vara de mirakel som lyser upp dystra naturkatastrofer .
I lördags räddades en liten pojke från en kloak .
I söndags räddade räddningsarbetarna en kvinna som varit fast under bråte i två dagar med sin mammas kropp bredvid sig .
Gendon Subandono , Indonesiens nationella skärmflygningslags tränare , hade tränat två av de saknade skärmflygarna inför Asiatiska spelen , som avslutades i Indonesien tidigare i månaden .
Andra som var fast på Roa Roa Hotel , inklusive mr Mandagi , var hans studenter .
" Som skärmflygningsveteran har jag en egen känslosam börda " , sa han .
Mr Gendon berättade att timmarna efter att skärmflygarna hörde att Roa Roa Hotel hade kollapsat skickade han desperat WhatsApp @-@ meddelanden till Palu @-@ deltagarna som deltog i strandfestivalen .
Men hans meddelanden fick bara en grå bock , i stället för två blå .
" Jag tror att det betyder att meddelandena inte levererades " , sa han .
Tjuvar tar $ 26.750 under bankomatpåfyllning vid Newport on the Levee
I fredags morse stal tjuvar $ 26.750 från en Brink ' s @-@ medarbetare som fyllde på en bankomat vid Newport on the Levee , enligt ett pressmeddelande från polisen i Newport .
Bilens förare hade tömt en bankomat i underhållningsanläggningen och skulle leverera mer pengar , sa kriminalare Dennis McCarthy i meddelandet .
Medan han var upptagen " sprang en annan man upp bakom Brink ' s @-@ medarbetaren " och stal en påse med pengar som skulle levereras .
Vittnen såg flera misstänkta fly från platsen , enligt pressmeddelandet , men polisen angav inte hur många som var inblandade i incidenten .
Alla som har information om förövarnas identitet ska kontakta polisen i Newport på 859 @-@ 292 @-@ 3680 .
Kanye West : Rapparen byter namn till Ye
Rapparen Kanye West byter namn - till Ye .
Han meddelade namnbytet på Twitter i lördags och sa : " Varelsen som formellt är känd som Kanye West " .
West , 41 , har kallats Ye under en längre tid och använde smeknamnet som titel för sitt åttonde album , som släpptes i juni .
Namnbytet kommer innan hans medverkan i Saturday Night Live , där han väntas lansera sitt nya album Yandhi .
Han ersätter sångaren Ariana Grande i programmet , som ställde in av " känslomässiga skäl " enligt programmets skapare .
Ye är en förkortning av Wests nuvarande professionella namn , men han har även sagt att ordet har en religiös betydelse för honom .
" Jag tror att " ye " är det ord som används mest i Bibeln , och i Bibeln betyder det " du " " , sa West tidigare i år när han pratade om titeln på sitt album med radiovärden Big Boy .
" Så jag är du , jag är vi , det är vi .
Det gick från Kanye , som betyder " den enda " , till bara Ye - en spegling av vårt goda , vårt onda , vårt förvirrade , allt .
Albumet är som en spegling av de vi är " .
Han är en av en rad kända rappare som har bytt namn .
Sean Combs har tidigare kallats Puff Daddy , P. Diddy och Diddy , men i år tillkännagav han att han föredrar att kallas Love och Brother Love .
JAY @-@ Z , som tidigare samarbetat med West , har tidigare skrivit sitt namn med och utan bindestreck och versaler .
Mexikos AMLO svär att inte använda militären mot civila
Mexikos nyligen valde president Andres Manuel Lopez Obrador har lovat att aldrig använda militären mot civilpersoner nu när landet närmar sig 50 @-@ årsdagen av en blodig vedergällning mot studenter .
Lopez Obrador lovade på Tlatelolco Plaza i lördags att " aldrig använda militären för att förtrycka det mexikanska folket " .
Trupper avfyrade vapen mot en fridfull demonstration på torget den andra oktober 1968 och dödade upp till 600 personer under en era då vänsterriktade studentrörelser slog rot i Latinamerika .
Lopez Obrador har svurit att stödja unga mexikaner med månatliga bidrag till studenter och genom att öppna fler kostnadsfria offentliga universitet .
Han har sagt att arbetslöshet och bristfälliga utbildningsmöjligheter lockar ungdomar till kriminella gäng .
USA borde fördubbla AI @-@ finansiering
Nu när Kina blir mer aktivt inom artificiell intelligens bör USA fördubbla den summa de spenderar på forskning inom fältet , enligt uppfinnaren och AI @-@ användaren Kai @-@ Fu Lee , som har arbetat för Google , Microsoft och Apple .
Kommentaren kommer efter att flera delar av USA:s regering har gjort uttalanden om AI , trots att USA inte har en övergripande formell AI @-@ strategi .
Kina presenterade sin plan i fjol med målet att bli ledande inom AI @-@ innovation innan 2030 .
" Det vore en bra början att fördubbla budgeten för AI @-@ forskning , med tanke på att alla andra länder ligger så långt bakom USA och vi letar efter nästa genombrott inom AI " , sa Lee .
En dubbelt så stor budget kan fördubbla chansen att nästa stora AI @-@ genombrott görs i USA , sa Lee till CNBC i en intervju tidigare i veckan .
Lee , vars bok " AI Superpowers : China , Silicon Valley and the New World Order " publicerades tidigare i månaden av Houghton Mifflin Harcourt , är VD för Sinovation Ventures , som har investerat i ett av Kinas mest framstående AI @-@ företag - Face + + .
På Carnegie Mellon University på 1980 @-@ talet arbetade han på ett AI @-@ system som slog den högst rankade amerikanska Othello @-@ spelaren , och senare satt han i ledningen för Microsoft Research och var VD för Googles Kina @-@ avdelning .
Lee nämnde tidigare teknologitävlingar från USA:s regering , som Robot Challenge från Advanced Research Projects Agency , och frågade vad nästa skulle bli för att kunna identifiera kommande visionärer .
I USA måste forskare ofta arbeta hårt för att få anslag från regeringen , sa Lee .
" Det är inte Kina som tar de akademiska ledarna från oss , utan företagen " , sa Lee .
De senaste åren har Facebook , Google och andra teknikföretag anställt ledande personligheter från universitet för att arbeta på AI .
Lee sa att nya immigrationspolicyer också kan hjälpa USA med AI @-@ innovationen .
" Jag tycker att green cards borde erbjudas automatiskt till doktorander inom AI " , sa han .
State Council i Kina utfärdade sin utvecklingsplan för nästa generation artificiell intelligens i juli 2017 .
I Kina ger National Natural Science Foundation anslag till personer på akademiska institutioner likt National Science Foundation och andra myndighetsorganisationer delar ut pengar till forskare i USA , men kvaliteten på det akademiska arbetet är lägre i Kina , sa Lee .
Tidigare i år etablerade USA:s försvarsdepartement ett Joint Artificial Intelligence Center som ska föra samman partner från industrin och den akademiska världen , och Vita huset meddelade bildandet av Select Committee on Artificial Intelligence .
Och tidigare denna månad tillkännagav DARPA en investering på $ 2 miljarder i ett initiativ de kallar AI Next .
NSF investerar för närvarande över $ 100 miljoner om året i AI @-@ forskning .
Amerikansk lagstiftning som skulle skapa en National Security Commission om artificiell intelligens har inte gjort några framsteg på flera månader .
Makedoniens folkomröstning om namnbyte
Makedoniens befolkning röstade i söndags i en folkomröstning om ifall landets namn ska ändras till " Republiken Nordmakedonien " , vilket skulle lösa en flera årtionden gammal dispyt med Grekland som har hindrat landets försök att gå med i Europeiska unionen och NATO .
Grekland har en provins som heter Makedonien och hävdar att namnet på dess granne i norr utgör ett krav på dess territorium och har därför hindrat Makedonien från att gå med i NATO och EU .
De två regeringarna slöt ett avtal i juni baserat på det föreslagna nya namnet , men nationalistiska motståndare hävdar att namnbytet skulle underminera Makedoniens slaviska majoritets identitet .
President Gjorge Ivanov har sagt att han inte tänker rösta i folkomröstningen och en bojkottkampanj har lett till tvivel om ifall minimideltagandet på 50 procent som krävs för att folkomröstningen ska anses vara giltig kommer att nås .
Frågan på valsedeln i folkomröstningen är följande : " Är du för medlemskap i NATO och EU med godkännande av avtalet med Grekland ? "
Men namnbytets anhängare , inklusive premiärminister Zoran Zaev , hävdar att det är värt att byta namn om det gör så att Makedonien , ett av länderna som bildades när Jugoslavien splittrades , kan gå med i EU och NATO .
" Jag är här för att rösta för vårt lands framtid , för ungdomar i Makedonien så att de kan leva fritt under Europeiska unionens paraply , för det innebär tryggare liv för oss alla " , sa Olivera Georgijevska , 79 , i Skopje .
Folkomröstningen är inte bindande , men tillräckligt med medlemmar i parlamentet har sagt att de tänker följa resultatet för att den ska anses avgörande .
Namnbytet kräver en majoritet på två tredjedelar av parlamentet .
Enligt den statliga valkommissionen hade inga oegentligheter rapporterats klockan 13 .
Men deltagandet var endast 16 procent , jämfört med 34 procent i det senaste parlamentsvalet 2016 då 66 procent av registrerade väljare röstade .
" Jag röstar för mina barns skull , vi hör hemma i Europa " , sa Gjose Tanevski , 62 , som röstade i huvudstaden Skopje .
Makedoniens premiärminister Zoran Zaev , hans fru Zorica och hans son Dushko röstar i folkomröstningen i Makedonien om landets namnbyte , som skulle öppna vägen för medlemskap i NATO och Europeiska unionen , i Strumica , Makedonien 30 september 2018 .
Utanför parlamentet i Skopje anordnade Vladimir Kavardarkov , 54 , en liten scen och ställe ut stolar framför tälten som har satts upp av de som bojkottar folkomröstningen .
" Vi är för NATO och EU , men vi vill gå med med huvudet i luften , inte smyga in genom bakdörren " , sa Kavardarkov .
" Vi är ett fattigt land , men vi har vår värdighet .
Om de inte välkomnar oss som Makedonien kan vi vända oss till andra , som Kina och Ryssland , och bli en del av en euro @-@ asiatisk integration " .
Enligt premiärminister Zaev skulle ett medlemskap i NATO leda till välbehövliga investeringar i Makedonien , som har en arbetslöshet på över 20 procent .
" Jag tror att den absoluta majoriteten kommer att rösta ja , för över 80 procent av våra invånare är för EU och NATO " , sa Zaev när han röstade .
Han sa att ett " Ja " -resultat vore en " bekräftelse på vår framtid " .
Enligt en undersökning som publicerades i måndags av Makedoniens institut för policyundersökning tänkte mellan 30 och 43 procent av väljare rösta i folkomröstningen , vilket faller under minimideltagandet som krävs .
Enligt en annan undersökning som utfördes av Telma TV i Makedonien tänkte 57 procent av deltagarna rösta på söndagen .
70 procent av dem tänkte rösta ja .
För att folkomröstningen ska räknas måste 50 procent av registrerade väljare plus en rösta .
Om folkomröstningen misslyckas blir det det första allvarliga bakslaget för den västerländskt inriktade regeringens policy sedan den tog över i maj i fjol .
Titta på : Manchester Citys Sergio Aguero tar sig genom hela Brightons försvar för att göra mål
Sergio Aguero och Raheem Sterling slog Brightons förslag i Manchester Citys vinst på 2 @-@ 0 på Etihad Stadium i Manchester , England i lördags .
Aguero fick det att se löjligt enkelt ut när han gjorde mål i 65:e minuten .
Den argentinska strikern fick en pass från mittfältet i början av sekvensen .
Han sprang mellan Brightons tre försvarare och gav sig ut på det öppna fältet .
Aguero var omgiven av fyra gröna tröjor .
Han tog sig runt en försvarare och sprang ifrån flera andra vid kanten av Brightons målområde .
Sedan pushade han en passning till Sterling till vänster .
Den engelska forwarden använde sin första spark i målområdet för att ge tillbaka bollen till Aguero , som använde högerfoten för att slå Brightons målvakt Mathew Ryan med ett skott i den högra sidan av nätet .
" Aguero har problem med fötterna " , sa Citys manager Pep Guardiola till journalisterna .
" Vi pratade om att han skulle spela i 55 @-@ 60 minuter .
Det är vad som hände .
Vi hade tur att han gjorde mål i det ögonblicket " .
Men det var Sterling som gav Sky Blues det inledande övertaget i Premier League @-@ kampen .
Målet kom i den 29:e minuten .
Aguero fick bollen djupt inne i Brightons revir på det spelet .
Han skickade iväg en fin spark längs den vänstra sidan till Leroy Sane .
Sane tog ett par sparkar och ledde Sterling till den bortre stolpen .
Sky Blues forward sparkade in bollen i nätet ögonblicket innan den hamnade utom räckhåll .
City möter Hoffenheim i gruppspelet i Champions League på Rhein @-@ Neckar @-@ Arena i Sinsheim , Tyskland klockan 12 : 55 på tisdag .
Scherzer vill spela mot Rockies
Nationals har eliminerats från slutspelet , så det fanns ingen anledning att tvinga fram en till start .
Men tävlingsinriktade Scherzer vill kasta på söndag mot Colorado Rockies , men bara om Rockies , som ligger en match före Los Angeles Dodgers i NL West , fortfarande har en chans till slutspelet .
Rockies fick en wild card @-@ plats med en vinst på 5 @-@ 2 över Nationals i fredags kväll , men är fortfarande ute efter sin första divisionstitel .
" Vi spelar om inget , men vi kan få en chans att gnugga gummit i vetskap om atmosfären här i Denver med publiken och att det andra laget skulle spela på högre nivå än något annat lag jag skulle möta i år .
Varför skulle jag inte vilja vara där ? "
Nationals har inte meddelat sin starter för söndag än , men enligt rapporter lutar de mot att låta Scherzer kasta under omständigheterna .
Scherzer , som skulle göra sin 34:e start , värmde upp i bullpenen i torsdags och skulle kasta på sin normala vilosöndag .
Washingtons högerhänta kastare är 18 @-@ 7 med 2,53 ERA och 300 strikeouts i 200 2 / 3 innings den här säsongen .
Trump håller tal i West Virginia
Presidenten hänvisade indirekt till situationen kring Brett Kavanaugh , som är nominerad till högsta domstolen , när han pratade om hur viktigt det är att republikaner röstar i de kommande midterm elections .
" Allt det vi har gjort står på spel i november .
Vi är fem veckor från ett av våra livs viktigaste val .
Det här är en av de stora , stora ... Jag kandiderar inte , men jag kandiderar . Det är därför jag åker runt och kämpar för suveräna kandidater " , sa han .
Trump fortsatte : " Ni ser en hemsk , hemsk grupp radikala demokrater , ni ser det hända här och nu .
De är fast beslutna att ta tillbaka makten vad som än krävs , ni ser deras elakhet , hemskhet .
De struntar i vem de måste såra , vem de måste köra över för att ta över makten och kontrollen . Det är det de vill ha , makt och kontroll . Vi ska inte låta dem få den " .
Demokrater , sa han , kämpar för att " stå emot och hindra " .
" Det har ni sett de senaste fyra dagarna " , sa han och kallade demokraterna " arga och elaka och hemska och falska " .
Han nämnde den demokratiska senatorn Dianne Feinstein , som sitter i Senate Judiciary Committee , vilket bemöttes av högt buande från åskådarna .
" Minns ni vad hon sa ?
" Läckte du dokumentet ? "
" Eh , eh , va ?
Nej , ej , nej , jag väntar en " ... Det var riktigt dåligt kroppsspråk , något av det värsta kroppsspråk jag har sett " .
Labour är inte längre en bred kyrka .
De tolererar inte personer som säger vad de tycker .
När Momentum @-@ aktivister i mitt lokala parti röstade för att censurera mig blev jag knappast förvånad .
Jag är ju trots allt den senaste i en rad MP från Labour som får höra att vi inte är välkomna , bara för att vi säger vad vi tycker .
Min kollega i parlamentet Joan Ryan behandlades på ett liknande sätt när hon stod på sig mot antisemitism .
I mitt fall kritiserades jag för att inte hålla med Jeremy Corbyn .
Om vikten av en ansvarsfull ekonomisk policy , om nationens säkerhet , om Europa - ironiskt nog liknande ämnen som Jeremy kritiserade tidigare ledare för .
I meddelandet om mötet med Nottingham East Labour i fredags stod det att " vi vill att mötena ska vara välkomnande och produktiva " .
Under större delen av mina åtta år som Labours lokala MP har GC @-@ mötena på fredagar varit precis det .
Men nu är tyvärr många möten inte det , och löftet om " vänligare , varsammare " politik har glömts bort för länge sedan , om det någonsin ens började .
Det har blivit alltmer uppenbart att avvikande åsikter inte tolereras inom Labour , och varje åsikt döms utifrån om partiets ledare accepterar den .
Detta började strax efter att Jeremy blev ledare , då kollegor som jag tidigare trodde hade en liknande politisk syn som jag väntade sig att jag skulle göra en helomvändning och ta ställningar som jag annars aldrig skulle ha hållit med om - vare sig det gällde nationens säkerhet eller EU:s inre marknad .
Varje gång jag talar offentligt - och det spelar egentligen ingen roll vad jag säger - följer en tirad av ovett på sociala medier som kräver att jag ska avsättas , kritiserar mittpolitiken och säger att jag inte ens borde vara med i Labour .
Och det här drabbar inte bara mig .
Faktum är att jag har mer tur än vissa av mina kollegor eftersom kommentarerna som riktas mot mig för det mesta är politiska .
Jag beundrar dessa kollegors professionalitet och beslutsamhet när de ställs inför en ström av sexistiska och rasistiska förolämpningar varenda dag men aldrig ger upp .
En av de största besvikelserna med denna eras politik är den nivå av förolämpningar som nu anses normal .
Jeremy Corbyn hävdade förra veckan att Labour ska främja en kultur av tolerans .
Men i verkligheten är vi inte längre denna breda kyrka och med varje misstroendeyrkande och förändring av urvalsreglerna blir partiet allt snävare .
Jag har fått många råd under de senaste två åren om att flyga under radarn och inte vara för rättfram , så " ordnar det sig " .
Men det var inte därför jag blev politiker .
Ända sedan jag gick med i Labour som skolelev för 32 år sedan , provocerad av Thatchers regerings försummelse som bokstavligt talat fick min grundskolas klassrum att falla samman , har jag försökt kämpa för bättre offentliga tjänster för de som behöver det mest - både på lokal nivå och som regeringsminister .
Jag har aldrig dolt mina politiska åsikter , och det inkluderar det senaste valet .
Ingen i Nottingham East kan på något sätt ha blivit förvirrad över mina åsikter om policyer och ämnen där jag inte håller med det nuvarande ledarskapet .
Till er som främjade yrkandet i fredags vill jag bara säga att när landet går mot ett Brexit som kommer att skada hushåll , verksamheter och offentliga tjänster förstår jag inte varför någon skulle vilja slösa tid och energi på min lojalitet mot Labours partiledare .
Men mitt främsta budskap är inte till Nottingham Momentum , utan till min valkrets - såväl Labour @-@ medlemmar som andra : Jag är stolt över att tjäna er och jag lovar att ingen mängd hot om att avsätta mig eller politisk bekvämlighet kommer att hindra mig från att göra det jag anser är bäst för er alla .
Chris Leslie är MP för Nottingham East
Ayr 38 @-@ 17 Melrose : Oslagna Ayr på topp
Två försök i sista minuten kan ha förvrängt resultatet en aning , men det finns inga tvivel om att Ayr förtjänade att triumfera i denna härligt underhållande Tennent ' s Premiership @-@ match .
De är nu på topp , den enda oslagna sidan av de tio .
I slutändan var det deras överlägsna försvar , såväl som deras förmåga att ta chanser , som gav hemmalaget vinsten , och tränaren Peter Murchie har all rätt att vara nöjd .
" Vi har testats under våra matcher hittills och är fortfarande oslagna , så vi är så klart glada " , sa han .
Robyn Christie från Melrose sa : " Ayr förtjänar det , de tog bättre chanser än vi " .
Grant Andersons försök i 14:e minuten , som konverterades av Frazier Climo , gav Ayr ledningen men ett gult kort för Skottlands kapten Rory Hughes , som släppts in av Warriors för matchen , lät Melrose låta siffrorna tala och Jason Baggot gjorde ett okonverterat försök .
Climo utökade Ayrs ledning med en straff , och i slutet av första halvleken gjorde han poäng och konverterade ett soloförsök för att ge Ayr en ledning på 17 @-@ 5 i pausen .
Men Melrose fick en bra start på andra halvleken och Patrick Andersons försök , som konverterades av Baggot , minskade ledningen till fem poäng .
Det blev sedan en lång väntan efter en allvarlig skada för Ruaridh Knott , som bars av planen , och efter omstarten ökade Ayr ledningen igen med ett försök från Stafford McDowall , som konverterades av Climo .
Ayrs agerande kapten Blair MacPherson fick sedan ett gult kort , och Melrose tvingade återigen den extra mannen att betala med ett okonverterat försök från Bruce Colvine , i slutet av en period med häftigt tryck .
Men hemmalaget återhämtade sig och när Struan Hutchinson fick ett gult kort för att ha tacklat Climo utan bollen gjorde McPherson en touch down från straff @-@ line @-@ outen bakom Ayrs maul .
Climo konverterade , vilket han gjorde igen nästan direkt efter omstarten , efter att Kyle Rowe samlade David Armstrongs box kick och skickade iväg flankern Gregor Henry för hemmalagets femte försök .
Still Game @-@ stjärna verkar redo för ny karriär i restaurangbranschen
Still Game @-@ stjärnan Ford Kiernan verkar redo att ge sig in i restaurangbranschen efter att det upptäckts att han har angetts som VD för en licensierad restaurangverksamhet .
56 @-@ åringen spelar Jack Jarvis i BBC:s populära serie , som han skriver och spelar i tillsammans med sin långvariga komedipartner Greg Hemphill .
Duon har tillkännagett att den kommande nionde säsongen blir seriens sista , och Kiernan verkar planera inför livet efter Craiglang .
Enligt officiella register är han VD för Adriftmorn Limited .
Skådespelaren nekade att kommentera , men en källa på Scottish Sun antydde att Kiernan ville ge sig in i Glasgows " blomstrande restaurangbransch " .
" Havet tillhör oss " : Kustlösa Bolivia hoppas att domstolen öppnar vägen till Stilla havet igen
Sjömän patrullerar ett riggtäckt högkvarter för flottan i La Paz .
Offentliga byggnader har en havsblå flagga .
Flottans baser från Titicacasjön till Amazonas bär mottot : " Havet tillhör oss .
Det är vår plikt att återhämta det " .
I kustlösa Bolivia är minnet av kustlinjen som förlorades till Chile i en blodig resurskonflikt på 1800 @-@ talet fortfarande starkt - och det är även längtan efter att återigen segla på Stilla havet .
Detta hopp är högre än på flera årtionden nu när Bolivia inväntar ett beslut från den internationella domstolen den första oktober , efter fem års övervägande .
" Bolivia har driften , en stämning av enhet och frid , och inväntar så klart resultatet med en positiv attityd " , sa Roberto Calzadilla , en boliviansk diplomat .
Många bolivianer kommer att se den internationella domstolens beslut på stora skärmar landet över , i hopp om att domstolen i Haag kommer att döma till fördel för Bolivias krav att Chile , efter åratal av oregelbundna diskussioner , måste förhandla med Bolivia om att tillåta dem ett eget utlopp till havet .
Måndagens beslut har även stor vikt för Evo Morales , Bolivias karismatiska infödda president som står inför en kontroversiell kamp för omval nästa år .
" Vi är väldigt nära att återvända till Stilla havet " , lovade han i slutet av augusti .
Men vissa analytiker anser att det är otroligt att domstolen dömer till Bolivias fördel , och att inte mycket skulle ändras även om den gör det .
FN:s domstol , med bas i Nederländerna , har inte rätt att tilldela chilenskt territorium och har stipulerat att den inte kommer att fastställa resultatet av möjliga diskussioner .
Det faktum att beslutet tillkännages endast sex månader efter de slutliga argumenten tyder på att fallet " inte var komplicerat " , sa Paz Zárate , en chilensk expert på internationell lag .
Och de senaste fyra åren kan snarare ha skadat än främjat Bolivias chanser .
" Frågan om åtkomst till havet har kapats av den nuvarande bolivianska administrationen " , sa Zárate .
Hon hävdar att Morales aggressiva retorik har tärt på Chiles kvarvarande välvilja .
Bolivia och Chile kommer så småningom att fortsätta diskussionen , men det blir extremt svårt att göra det efter detta .
De två länderna har inte utbytt ambassadörer sedan 1962 .
Före detta presidenten Eduardo Rodríguez Veltzé , Bolivias representant i Haag , ansåg inte att domstolens beslut hade fattats ovanligt snabbt .
Måndagen kommer att ge Bolivia " en enastående möjlighet att inleda en ny era för relationen med Chile " och en chans att " sätta stopp för 139 år av meningsskiljaktigheter med ömsesidiga fördelar " , sa han .
Calzadilla förnekade även att Morales - fortfarande en av Latinamerikas populäraste presidenter - använde frågan om havet som politisk krycka .
" Bolivia kommer aldrig att ge upp sin rätt att ha åtkomst till Stilla havet " , sa han .
" Beslutet är en chans att inse att vi måste gå vidare från det förflutna " .
Nordkorea säger att kärnvapennedrustning kräver tillit till USA
Nordkoreas utrikesminister Ri Yong Ho säger att nationen inte kommer att nedrusta sina kärnvapen först om de inte kan lita på Washington .
Ri talade till FN:s generalförsamling i lördags .
Han uppmanade USA att uppfylla de löften som gjordes under ett toppmöte i Singapore mellan de två rivaliserande ledarna .
Hans kommentarer kom då USA:s utrikesminister Mike Pompeo verkar vara på gränsen att lösa dödläget för kärnvapendiplomatin mer än tre månader efter mötet i Singapore med Nordkoreas ledare Kim Jong Un .
Ri säger att det är en " önskedröm " att fortsatta sanktioner och USA:s protester mot ett uttalande om att avsluta Koreakriget någonsin kommer att tämja Nordkorea .
Washington tvekar inför att gå med på uttalandet utan att Pyongyang först inleder betydande kärnvapennedrustning .
Både Kim och USA:s president Donald Trump vill ha ett till toppmöte .
Men det finns utbredd skepticism mot att Pyongyang verkligen tänker göra sig av med en vapenarsenal som landet troligen ser som sin enda chans att garantera sin säkerhet .
Pompeo planerar att besöka Pyongyang nästa månad för att förbereda inför att andra toppmöte mellan Kim och Trump .
Paris modevisningar avslöjar senaste linje enorma huvudbonader på väg till butiker nära dig
Om du vill förstora din hattsamling eller helt blockera solen har vi rätt grej för dig .
Designerna Valentino och Thom Browne har avslöjat ett utbud av knasiga , överdimensionerade huvudbonader för sin SS19 @-@ kollektion på catwalken , som bländade stilikonerna på Paris modevecka .
Otroligt opraktiska hattar har tagit över Instagram denna sommar , och designerna har skickat iväg sina iögonfallande skapelser på catwalken .
Valentinos främsta skapelse var en överdriven beige hatt med ett fjäderliknande brett hattbrätte som helt tog över modellernas huvuden .
Andra överdimensionerade accessoarer inkluderade juvelprydda vattenmeloner , en trollkarlshatt och till och med en ananas - men de är inte avsedda att hålla huvudet varmt .
Thom Browne avslöjade även ett urval bisarra maskar , i lagom tid för Halloween .
Många av de färgglada maskarna hade ihopsydda läppar och liknade snarare Hannibal Lecter än haute couture .
En skapelse liknade en våtdräkt med snorkel och dykmask , och en annan såg ut som en smält glasstrut .
Och om du fortsätter det enorma modet har du tur .
Modeexperter förutsäger att de enorma hättorna kan vara på väg till butiker nära dig .
De överdimensionerade hattarna kommer strax efter La Bomba - halmhatten med ett brätte på 60 cm som har setts på alla från Rihanna till Emily Ratajkowski .
Kultmärket som låg bakom den otroligt opraktiska hatten som har tagit över sociala medier skickade ut ännu en stor skapelse på catwalken - en halmstrandväska som var nästan lika stor som modellen i baddräkt som höll i den .
Raffiaväskan i terrakotta , med raffiafransar och ett vitt läderhandtag , utmärkte sig i Jacquemus La Riviera SS19 @-@ kollektion på Paris modevecka .
Kändisstylisten Luke Armitage sa till FEMAIL : " Jag väntar mig att se stora hattar och strandväskor i butikerna nästa sommar - designern har haft en så stor inverkan att det vore svårt att ignorera efterfrågan på överdimensionerade accessoarer " .
John Edward : Språkfärdigheter avgörande för globala medborgare
Skottlands oberoende skolor bibehåller enastående akademiska resultat och detta fortsatte 2018 med ännu en uppsättning enastående provresultat , som bara stärks av individuella och kollektiva framsteg inom sport , konst , musik och andra samhällsengagemang .
Med upp till 30.000 elever i Skottland strävar skolorna , som representeras av The Scottish Council of Independent Schools ( SCIS ) , efter att tillhandahålla bästa möjliga service för sina elever och deras föräldrar .
Oberoende skolor strävar efter att förbereda sina elever inför vidare utbildning , deras valda karriär och deras roll som globala medborgare .
Som en utbildningssektor som kan utforma och implementera anpassade läroplaner ser vi att moderna språk fortsätter vara populära och efterfrågade ämnen på skolorna .
Nelson Mandela sa : " Om du pratar med en man på ett språk han förstår går det till hans huvud .
Om du pratar med honom på hans eget språk går det till hans hjärta " .
Det är en mäktig påminnelse om att vi inte bara kan förlita oss på engelska när vi skapar relationer och tillit med personer från andra länder .
Detta års provresultat visar att språk ligger högst på listan , med högst antal godkända resultat inom oberoende skolor .
Sammanlagt 68 procent av elever som studerade främmande språk fick A i slutprovet Higher Grade .
Data , som samlades in från SCIS 74 medlemsskolor , visade att 72 procent av elever som studerade mandarin fick ett A i Higher Grade , och 72 procent av de som studerade tyska , 69 procent av de som studerade franska och 63 procent av de som studerade spanska fick också ett A.
Detta visar att oberoende skolor i Skottland stödjer främmande språk som avgörande färdigheter som barn och ungdomar utan tvekan kommer att behöva i framtiden .
Språk som ämnesval anses nu vara lika viktiga som naturkunskap , teknik , ingenjörskunskap och matematik på läroplaner i oberoende skolor och bortom .
En undersökning genomförd av Storbritanniens Commission for Employment and Skills 2014 kom fram till att arbetsgivare av olika anledningar hade svårt att fylla sina lediga tjänster , med 17 procent som tillskrevs en brist på färdigheter i språk .
Med detta sagt , blir språkfärdigheter all mer nödvändigt för att förbereda unga människor för deras framtida karriärer .
Med allt fler framtida arbetstillfällen som kräver språkfärdigheter , blir dessa kompetenser nödvändiga i en globaliserad värld .
Oavsett karriärvalet , kommer de att ha en verklig fördel i framtiden om de har anammat sig ett andraspråk .
Att kunna kommunicera direkt med människor från andra länder , ger automatiskt en flerspråkig person en konkurrensfördel .
Enligt en undersökning av fler än 4 000 vuxna britter publicerad av YouGov 2013 , svarade 75 procent att de inte kunde tala ett främmande språk bra nog för att hålla en konversation i det , och där franska var det enda språket som total kom upp i ett två @-@ siffrigt procenttal ( 15 procent ) .
Därför är det så viktigt att investera i språkundervisning för våra barn .
Att kunna tala flera språk , särskilt de som används i utvecklingsländer , ger ditt barn en bättre chans att hitta en meningsfull sysselsättning i framtiden .
I Skottland kommer varje skola lära ut olika kombinationer av språk .
Ett antal skolor kommer att fokusera på de mer klassiska moderna språken , medan andra kommer att undervisa i språk som anses vara viktigast för Storbritannien inför 2020 , till exempel kinesiska eller japanska .
Oavsett ditt barns intresse kommer det alltid att finnas ett antal språk att välja mellan inom fristående skolor , med lärare som är specialister på detta område .
Skotska självständiga skolor strävar efter att tillhandahålla en läromiljö som kommer att förbereda barn och få dem med de färdigheter som krävs för att lyckas , oavsett vad framtiden har på lut .
I en global ekonomisk miljö är det utan tvekan språk som fortsätter att vara avgörande för landets framtid , så det måste speglas i utbildningen .
I själva verket borde moderna språk verkligen betraktas som " internationell kommunikationsförmåga " .
Oberoende skolor kommer att fortsätta erbjuda detta val , mångfald och excellens för Skottlands ungdomar .
Il faut bien le faire .
John Edward är chef för Scottish Council of Independent Schools
LeBron gör Lakersdebut på söndag i San Diego
Väntan är nästan över för fans som ser fram emot att se LeBron James göra debut för Los Angeles Lakers .
Lakers tränare Luke Walton har meddelat att James kommer att spela i söndagens första säsongsmatch mot Denver Nuggets i San Diego .
Men hur många minuter han spelar har ännu inte bestämts .
" Det kommer att bli mer än en och mindre än 48 " , sa Walton på Lakers officiella hemsida .
Lakers reporter Mike Trudell tweetade att James sannolikt kommer att spela ett begränsat antal minuter .
Efter att ha tränat tidigare i veckan blev James tillfrågad om sina planer för Lakers " försäsongsschema .
" Jag behöver inte försäsongsspel i detta stadie av min karriär för att bli redo " , sa han .
Trumps West Virginia kampanjevenemang , YouTube @-@ kanal
President Donald Trump gör sitt första kampanjevenemang ikväll i Wheeling , West Virginia .
Det är Trumps första av fem planerade uppträdanden under nästa vecka , inklusive evenemang på platser han har stort stöd , såsom Tennessee och Mississippi .
I väntan på en bekräftande omröstning av sin kandidat till högsta domstolens lediga post , syftar Trump till att bygga upp stöd för kommande mellanårsval , eftersom republikanerna riskerar att förlora kontrollen över kongressen inför det stundande valet i november .
Vilken tid är Trumps West Virginia rally i kväll och hur kan du titta på det på nätet ?
Trumps Wheeling , West Virginia kampanjevenemang är planerat till 19 : 00 , ikväll lördag , 29 september 2018 .
Du kan titta på Trumps West Virginia @-@ rally online nedan via live stream på YouTube .
Trump kommer sannolikt att ta itu med denna veckas förhör av kandidaten till högsta domstolen Brett Kavanaugh , som blev spända efter beskyllningar om hans sexuella övergrepp , med en förväntad försening av omröstningen från senaten på upp till en vecka medan FBI:s utredning av fallet pågår .
Men det primära syftet med dessa evenemang är att hjälpa republikanerna att få lite kött på benen inför novembervalet .
Således sade president Trump att dessa fem sammankomster i nästa vecka syftar till att " engagera volontärer och anhängare då republikanerna försöker skydda och utöka majoriteten i senaten och representanthuset " , enligt Reuters .
" Kontroll av kongressen är så viktig för hans agenda att presidenten kommer att resa till så många stater som möjligt när vi går in i den hektiska kampanjperioden " , sa en talesman för Trump @-@ kampanjen som inte ville bli namngiven till Reuters .
Nattens evenemang , schemalagt på Wesbanco Arena i Wheeling , kan dra in fans från " Ohio och Pennsylvania och locka till sig uppmärksamhet från Pittsburghs media " , enligt West Virginia Metro News .
Lördag blir andra gången under den senaste månaden som Trump har besökt West Virginia , staten där han vann med mer än 40 procentenheter år 2016 .
Trump försöker hjälpa den republikanska senatkandidaten för West Virginia , Patrick Morrisey , som har halkat efter i opinionsundersökningarna .
" Det är inte ett gott tecken för Morrisey att presidenten måste komma dit för att försöka ge honom en ökning i opinionsundersökningarna " , säger Simon Haeder , en statsvetare vid West Virginia University , enligt Reuters .
Ryder Cup 2018 : Team USA kämpar för att hålla förhoppningarna vid liv inför söndagens singlar
Efter tre ensidiga sessioner kunde partävlingarna i lördags eftermiddag ha varit vad som krävdes för denna Ryder Cup .
Momentets svängande pendel är ett helt uppfunnet sportkoncept , men något som spelarna verkligen tror på , och mer än någonsin inför tävlingar som dessa .
Så vilket momentum handlar det om nu ?
" De hade en sexpoängsledning och nu är det fyra , så vi bär det som ett litet momentum gissar jag " sa Jordan Spieth när han avslutat för dagen .
Europa har fördelen , naturligtvis , fyra poängs förskott med tolv mer att vinna .
Amerikanerna , som Spieth säger , känner att de har lite vind i seglen , men de har mycket att uppmuntras av , inte minst i form av Spieth och Justin Thomas som spelade tillsammans hela dagen och kammade hem tre poäng av fyra var .
Spieth har varit vass från tee till green och föregår med gott exempel .
Vinstropen skallade än högre när hans runda fortsatte och han sänkte en avgörande putt för att ta matchen fyra all @-@ square när han och Thomas hade legat efter med två efter två spel .
Hans putt som vann dem matchen på 15 möttes med ett liknande vrål , med övertygelsen om att det amerikanska laget ännu inte är ute ur spelet .
" Du måste verkligen gräva djupt och oroa dig för din egen match " , sa Spieth .
Det är allt som alla dessa spelare har kvar nu .
18 hål till seger .
De enda spelarna med fler poäng än Spieth och Thomas under de senaste två dagarna är Francesco Molinari och Tommy Fleetwood , Ryder Cups obestridliga berättelse .
Europas udda men bedårande par är fyra från fyra och nu kan inget gå fel .
" Moliwood " var det enda paret som inte gjorde en bogey på lördag eftermiddag och de undvek också bogeys på lördag morgon , fredag eftermiddag och back nine på fredagsmorgonen .
Dessa prestationer och publikens reaktioner slår fast att de är spelarna att slå på söndag och det finns ingen mer populär spelare som skulle kunna kamma hem en potentiell europeisk seger när solen går ner över Le Golf National än Fleetwood eller Molinari .
Företrädesvis båda , samtidigt på olika hål .
Det är dock för tidigt att tala om europeisk seger .
Bubba Watson och Webb Simpson gjorde processen kort med Sergio Garcia , morgonens fyrbolls @-@ hjälte , tillsammans med Alex Noren .
En bogey och två dubblar på front nio sänkte spanjoren och svensken i ett hål som de aldrig ens kom i närheten att kravla sig ur .
På söndag finns det emellertid ingen som hjälper dig ut ur hålet .
Fyrboll och foursome är så fascinerande att se på nära håll på grund av samspelet mellan paren , de råd de ger , de råd de inte ger och hur en strategi kan förändras på ett ögonblick .
Europa har spelat bättre som lag hittills och tagit en betydande ledning inför sista dagen men denna foursomesession visade också att Team USA har en kämpaglöd som vissa , särskilt på USA:s sida , hade tvivlat på .
Europa tar ledningen med 10 @-@ 6 i Ryder Cup sista dagen
Europa kommer att ha en stark fördel på Ryder Cups sista dag efter att ha kommit ut från lördagens fyrboll och foursomes matchad med en 10 @-@ 6 @-@ ledning över USA .
Den inspirerade duon Tommy Fleetwood och Francesco Molinari ledde med två segrar över en belägrad Tiger Woods och kammade hem hela fyra poäng vid Le Golf National .
Thomas Bjorns europeiska lag , som kämpade för att behålla pokalen som de förlorade vid Hazeltine för två år sedan dominerade ett amerikanskt lag som aldrig riktigt kom igång under morgonens fyrboll med 3 @-@ 1 .
USA erbjöd mer motstånd i foursomen och vann två matcher , men det räckte inte för seger .
Jim Furyks lag behöver åtta poäng från söndagens 12 singelmatcher för att behålla pokalen .
Fleetwood är den första europeiska nybörjaren att vinna fyra poäng i rad medan han och Molinari , döpta till " Molliwood " , efter en sensationell helg är bara det andra paret att vinna fyra poäng från deras första fyra matcher i Ryder Cups historia .
Efter att ha krossat Woods och Patrick Reed i fyrboll , slog de en utmattad Woods och American rookie Bryson Dechambeau med en ännu mer eftertrycklig 5 & 4 .
Woods , som slog sig igenom två matcher på lördag , visade prov på enstaka stunder av briljans , men han har nu förlorat 19 av sina 29 matcher i fyrboll och foursome , och därav sju i rad .
Justin Rose , vilade under morgonens fyrboll och återvände till partnern Henrik Stenson i foursomes till ett 2 & 1 @-@ seger över Dustin Johnson och Brooks Koepka - rankad etta och trea i världen .
Europa hade inte medvind hela vägen , men det var en trevlig , blåsig dag strax sydväst om Paris .
Trefaldige vinnaren Jordan Spieth och Justin Thomas satte riktmärket för amerikanerna med två poäng på lördag .
De kammade hem segern med 2 & 1 över Spaniens Jon Rahm och Ian Poulter i fyrboll och återvände senare för att slå Poulter och Rory McIlroy 4 & 3 i foursome efter att ha förlorat de två öppningshålen .
Endast två gånger i Ryder Cups historia har ett lag kommit tillbaka från ett underläge på fyra poäng i singelmatcherna , dock behöver Furyks sida bara ett oavgjort resultat för att behålla pokalen .
Efter att ha varit näst bäst i två dagar ser det ut som en motattack på söndagen kan bli svår att få igenom .
Nordkorea säger att de " aldrig " kommer att avväpna ensidigt utan förtroende
Nordkoreas utrikesminister berättade för Förenta nationerna i lördags att fortsatta sanktioner fördjupade deras misstro gentemot USA och det inte var möjligt att landet skulle ge upp sina kärnvapen ensidigt under sådana omständigheter .
Ri Yong Ho berättade för världsorganisationens årliga generalförsamling att Nordkorea under det senaste året hade vidtagit " betydande åtgärder för att visa sin välvilja " , till exempel genom att stoppa kärnvapen- och missilprov , demontera installationerna för kärnvapenprov och lova att inte sprida kärnvapen och kärnvapenteknik .
" Vi ser emellertid inte något motsvarande svar från USA " , sa han .
" Utan något förtroende för USA kommer det inte att finnas något förtroende för vår nationella säkerhet och under sådana omständigheter finns det inte en chans att vi ensidigt avväpnar oss själva först " .
Medan Ri upprepade välbekanta nordkoreanska klagomål om Washingtons motstånd mot ett tillvägagångssätt uppdelat i etapper för den kärnkraft som skulle leda till att Nordkorea skulle belönas då det tog gradvisa steg , verkade hans uttalande betydelsefullt , eftersom det inte avvisade en ensidig kärnvapenlösning helt såsom Pyongyang tidigare gjort .
Ri hänvisade till ett gemensamt uttalande utfärdat av Kim Jong Un och Donald Trump vid det första toppmötet mellan en sittande amerikansk president och en nordkoreansk ledare i Singapore 12 juni , där Kim lovade att arbeta mot " avveckling av kärnvapen på den koreanska halvön " medan Trump lovade garantier för Nordkoreas säkerhet .
Nordkorea har sökt ett formellt slut på Korea @-@ kriget 1950 @-@ 53 , men USA har sagt att Pyongyang först måste avveckla sina kärnvapen .
Washington har också tackat nej till förhandlingar om att lätta på hårda internationella sanktioner mot Nordkorea .
" USA insisterar på " avveckling först " och ökar trycket genom sanktioner för att uppnå sitt syfte genom tvång och invänder till och med mot " deklarationen om att avsluta kriget " " , säger Ri .
" Uppfattningen om att sanktioner kan få oss på knäna är en önskedröm för de människor som saknar kunskap om oss .
Men problemet är att de fortsatta sanktionerna fördjupar vår misstro " .
Ri nämnde inte planer på ett andra toppmöte mellan Kim och Trump som USA:s ledare framhävde i FN tidigare under veckan .
Ministern pekade istället på tre möten mellan Kim och Sydkoreas ledare Moon Jae @-@ in under de senaste fem månaderna och tillade : " Om parten i denna fråga om kärnvapennedrustning varit Sydkorea och inte USA , skulle den koreanska halvöns kärnvapennedrustning inte ha kommit till ett sådant dödläge " .
Ändå var tonen i Ri:s tal dramatiskt annorlunda än förra året när han berättade för FN:s generalförsamling att Nordkoreas framtida förmåga att nå USA:s fastland med raketer var oundvikligt efter " Mr Evil President " Trump kallade Kim en " raketman " på ett självmordsuppdrag .
I år i Förenta nationerna , gav Trump , som i fjol hotade att " helt förstöra " Nordkorea , beröm till Kim för hans mod att vidta åtgärder för avväpning , men det sade att mycket arbete fortfarande återstår och att sanktioner måste kvarstå tills Nordkorea avväpnas .
På onsdagen sade Trump att han inte hade någon tidsram för detta och sade att " om det tar två år , tre år eller fem månader " , spelar ingen roll " .
Kina och Ryssland hävdar att FN:s Säkerhetsrådet bör belöna Pyongyang för de åtgärder som vidtagits .
USA:s Statssekreterare Mike Pompeo sa emellertid till FN:s säkerhetsråd på torsdagen att : " Upprätthållandet av säkerhetsrådets sanktioner måste fortsätta med kraft och utan att misslyckas tills vi förverkligar en fullständig , slutgiltig , verifierad nedrustning " .
Säkerhetsrådet har enhälligt förstärkt sanktionerna mot Nordkorea sedan 2006 i ett försök att kväva finansieringen av Pyongyangs kärnvapen- och ballistiska missilprogram .
Pompeo träffade Ri i samband med FN:s generalförsamling och sa därefter att han skulle besöka Pyongyang igen nästa månad för att förbereda sig för ett andra toppmöte .
Pompeo har besökt Nordkorea tre gånger redan i år , men hans sista resa gick inte bra .
Han lämnade Pyongyang i juli och sade att framsteg hade gjorts . Nordkorea anklagade honom dock några timmar senare för ställa " gangsterliknande krav " .
Nordkorea lovade ett möte med Moon denna månad för att demontera en missilanläggning och även ett kärnkrafkomplex om USA vidtog " motsvarande åtgärder " .
Han sa att Kim hade sagt till honom att de " motsvarande åtgärder " han sökte var säkerhetsgarantier som Trump lovade i Singapore och rör sig mot normalisering av relationerna med Washington .
Harvardstudenter tar kurs om att få tillräckligt med vila
En ny kurs på Harvard University i år har fått alla doktorander att förbättra sina sömnvanor i ett försök att bekämpa den växande machokulturen att studera genom koffeinfyllda " dygningar " .
En akademisk studie fann att studenter vid världens ledande universitet ofta är aningslösa när det gäller själva grunderna för hur man ska ta hand om sig .
Charles Czeisler , professor i sömnmedicin vid Harvard Medical School och en specialist på Brigham och Women ' s Hospital , utformade kursen , som han anser är den första i sitt slag i USA .
Han inspirerades att starta kursen efter att ha pratat om vilken inverkan sömnbrist hade på inlärning .
" I slutet av det kom en tjej upp till mig och sa : Varför får jag inte veta detta förrän nu , under mitt sista år ? "
Hon sa att ingen någonsin hade berättat för henne om vikten av sömn - vilket förvånade mig , berättade han för The Telegraph .
Kursen , som anordnades för första gången i år , förklarar för studenterna vikten av hur bra sömnvanor hjälper akademisk och atletisk prestation , samt förbättrar deras allmänna välbefinnande .
Paul Barreira , professor i psykiatri vid Harvard Medical School och verkställande direktör för universitetets hälsovårdstjänster , sa att universitetet bestämde sig för att introducera kursen efter att ha upptäckt att eleverna led av allvarlig sömnbrist under veckan .
Den timslånga kursen omfattar en rad interaktiva uppgifter .
I en del av kursen finns en bild av ett studentrum , där eleverna klickar på kaffekoppar , gardiner , tränare och böcker för att få veta om effekterna av koffein och ljus , hur atletisk prestation påverkas av sömnbrist och vikten av goda sömnvanor .
I en annan del får deltagarna veta hur långsiktig sömnbrist kan öka riskerna för hjärtattacker , stroke , depression och cancer .
En karta över campus , med interaktiva ikoner , uppmuntrar deltagarna att tänka på sin dagliga rutin .
" Vi vet att det inte kommer att förändra elevernas beteende direkt .
Men vi tror att de har rätt att veta - precis som man har rätt att veta om hälsoeffekterna av att välja att röka cigaretter " , tillade Professor Czeisler .
Stolthetskulturen i att " dygna " finns fortfarande , säger han och tillade att modern teknik och ständigt ökande tryck på eleverna betydde att sömnbrist var ett växande problem .
Att säkerställa att du har tillräckligt med sömn , av god kvalitet , borde vara studentens " hemliga vapen " för att bekämpa stress , utmattning och ångest , sade han - även för att undvika viktuppgång eftersom sömnlöshet sätter hjärnan i svältläge och gör dem ständigt hungriga .
Raymond So , en 19 @-@ årig kalifornier som studerar kemisk och fysisk biologi , hjälpte professor Czeisler att utforma kursen och har läst en av hans kurser förra året under sitt första år på Harvard .
Han sa att kursen var en ögonöppnare och inspirerat honom att kampanja för en campusövergripande kurs .
Han hoppas att nästa steg är att be alla doktorander att slutföra ett liknande studieprogram innan de påbörjar sina studier vid den högpresterande institutionen .
Professor Czeisler rekommenderade att eleverna överväger att sätta ett larm för när man ska lägga sig och när man ska vakna och vara medvetna om de skadliga effekterna av " blått ljus " som emitteras av elektroniska skärmar och LED @-@ belysning , som kan få dig att vända på dygnet , vilket leder till insomningsproblem .
Livingston 1 - 0 Rangers : Mengas mål sänker Gerrards män
Rangers led ännu en förlust i dag då Dolly Mengas strike skickade Steven Gerrards ojämna sida till ett 1 @-@ 0 @-@ nederlag i Livingston .
Ibrox @-@ sidan var ute efter att ta hem sin första seger på vägen sedan februaris 4 @-@ 1 @-@ triumf på St Johnstone , men Gary Holts lag levererade Gerrards andra nederlag i 18 matcher som manager för att lämna hans lag åtta poäng efter Ladbrokes Premiership @-@ ledaren Harts .
Menga slog till sju minuter före halvtid och Rangers lyckades aldrig jämna ut resultatet .
Medan Rangers nu faller ner till sjätte plats , klättrar Livingston till tredje och ligger bara bakom Hibernian på målskillnad .
Och det kan finnas fler problem på lut för Rangers efter att linjeman Calum Spence var tvungen att behandlas för ett huvudsår efter att ett föremål kastats från den bortre änden .
Gerrard gjorde åtta ändringar i semifinalen i Betfred Cup .
Holt å andra sidan gick med samma Livi 11 som tog en poäng av Hearts förra veckan och han skulle ha varit glad över sättet hans välsmorda spel överglänste motståndarna varje gång .
Rangers må ha dominerat , men Livingston gjorde mer med bollkontrollen de hade .
Det borde ha blivit mål redan två minuter in i matchen när Mengas första pass släppte igenom Scott Pittman till Allan McGregors mål , men mittfältaren missade sin stora chans och sköt utanför .
En frispark på djupet från Keaghan Jacobs nådde sedan lagkaptenen Craig Halkett , men hans defensiva partner Alan Lithgow nådde bara bakre stolpen .
Rangers tog kontroll över matchen , men det såg ut att vara mer hopp än tro i deras spel under matchens sista tredjedel .
Alfredo Morelo kände säkert att han borde ha haft straff när han och Steven Lawless kolliderade , men domaren Steven Thomson viftade bort colombianens uppmaning .
Rangers lyckades bara göra två mål i första halvlek men den före detta Ibroxmålvakten Liam Kelly tog lätt emot Lassana Coulibalys nick och en tam spark från Ovie Ejaria .
Livis öppningsskott i 34:e minuten må gått emot spelets anda , men ingen kan neka till att deras knegande förtjänade det .
Återigen misslyckades Rangers att hantera Jacobs fasta situation .
Scott Arfield reagerade inte när Declan Gallagher passade till Scott Robinson , som höll sig lugn och valde Menga för ett enkelt avslut .
Gerrard agerade vid pausen när han bytte Coulibaly till Ryan Kent och bytet gav nästan omedelbar effekt när yttern slog in bollen till Morelos , men den imponerande Kelly sprang från sin linje för att blockera försöket .
Men Livingston fortsatte att få motspelarna att spela exakt den typ av spel de tycker om , med Lithgow och Halkett som svepte upp lång passning efter lång passning .
Holts sida skulle kunna ha stärkt sin ledning i sista etappen , men McGregor klarade väl att hindra Jacobs innan Lithgow nickade utanför efter hörnan .
Rangers @-@ ersättaren Glenn Middleton hade ännu ett sent krav på straff när han tampades med Jacobs , men återigen tittade Thomson bort .
Almanac : Uppfinnaren av Geiger Counter
Och nu en sida från söndagens almanacka : 30 september 1882 , 136 år sedan idag ... dagen då den framtida fysikern Johannes Wilhelm " Hans " Geiger föddes i Tyskland .
Geiger utvecklade en metod för att detektera och mäta radioaktivitet , en uppfinning som så småningom ledde till manicken kallad Geigermätare .
Geigermätare har blivit en grundsten för vetenskapen sedan dess och figurerar även stort inom popkultur , liksom i 1950 @-@ filmen " Bells of Coronado " , med huvudrollen i de till synes osannolika cowpokeforskarna Roy Rogers och Dale Evans :
MAN " Vad i all världen är det där ? "
Rogers : " Det är en Geigermätare , som används för att lokalisera radioaktiva mineraler , som uran .
När du sätter på dig dessa hörlurar kan du faktiskt höra effekterna av atomerna som avges av radioaktiviteten i mineralerna . " Evans :
Evans : " Ja , det poppar nu ! "
" Hans " Geiger dog 1945 , bara några dagar innan sin 63 @-@ årsdag .
Men uppfinningen som bär hans namn lever vidare .
Nytt cancervaccin kan lära immunförsvaret att " se " cancerceller
Nytt cancervaccin kan lära immunförsvaret att " se " cancerceller och döda dem
Vaccin lär immunsystemet att känna igen cancerceller som en del av behandlingen
Metoden innebär att extrahera immunceller från en patient och modifiera dem i laboratoriet
De kan då " se " ett protein som är gemensamt för många cancerformer och sedan återinjiceras
Ett försöksvaccin visar lovande resultat hos patienter med olika cancerformer .
En kvinna behandlad med vaccinet , som lär immunsystemet att känna igen cancer , såg sina äggstockscancerceller försvinna i över 18 månader .
Metoden involverar att extrahera immunceller från en patient och modifiera dem i laboratoriet så att de kan " se " ett protein som är gemensamt för många cancerformer som kallas HER2 , och sedan återinjicera cellerna .
Professor Jay Berzofsky , från US National Cancer Institute i Bethesda , Maryland , sa : " Våra resultat tyder på att vi har ett mycket lovande vaccin " .
HER2 " främjar tillväxten av flera typer av cancer , inklusive bröst- , äggstocks- , lung- och tjocktarmscancer , förklarade Prof Berzofsky .
En liknande metod att ta immunceller från patienter och " lära " dem hur man riktar sig mot cancerceller har fungerat vid behandling av en typ av leukemi .
Kanye West stöttade Trump genom att bära en MAGA @-@ keps , efter sitt SNL @-@ framträdande .
Det gick inte så bra
Kanye West buades ut ur studion under Saturday Night Live efter ett svamlande framträdande där han lovordade USA:s President Donald Trump och sa att han själv skulle kandidera för posten 2020 .
Efter att ha utfört sin tredje låt för kvällen , kallad Ghost Town där han hade på sig en Make America Great @-@ keps , raljerade han emot demokraterna och upprepade sitt stöd för Trump .
" Så många gånger när jag pratar jag med en vit person säger de : " Hur kan du tycka om Trump , han är rasistisk ? "
Tja , om jag var bekymrad över rasism skulle jag ha flyttat från Amerika för länge sen , sa han .
SNL startade showen med en sketch med Matt Damon där Hollywoodstjärnan gjorde narr av Brett Kavanaughs vittnesbörd inför senatens rättsliga kommitté om de anklagelser om sexuella övergrepp som gjorts av Christine Blasey Ford .
Även om det inte sändes , laddades uppspelningen av Wests utläggning upp på sociala medier av komikern Chris Rock .
Det är oklart om Rock försökte driva med West med inlägget .
West hade också beklagat sig inför publiken att han hade blivit trakasserad backstage för sin huvudbonad .
" De mobbade mig backstage .
De sa : " Gå inte ut dit med den kepsen på " .
De mobbade mig !
Och sen säger de att jag sjunkit lågt " , sa han , enligt Washington Examinator .
West fortsatte : " Vill du också sjunka lågt ? " och sa att han skulle " sätta min supermancape på , för det betyder att du inte kan säga vad jag får göra . Vill du att världen ska gå framåt ?
Testa med kärlek " .
Hans kommentarer lockade fler burop åtminstone två gånger från publiken och medarbetare från SNL tycktes generade , rapporterade Variety . En person sa : " Det blev dödstyst i studion " .
West hade kommit in som en sen ersättare för sångaren Ariana Grande , vars före detta pojkvän , rapparen Mac Miller hade dött för några dagar sedan .
West förbryllade många med sitt framträdande av låten I Love it , utklädd till en Perrierflaska .
West fick stöd från chefen för konservativa gruppen TPUSA , Candace Turner som tweetade : " Till en av de modigaste själarna : TACK FÖR ATT DU STOD PÅ DIG MOT MOBBEN " .
Men pratshowens värd , Karen Hunter , tweetade att West helt enkelt " var sig själv och det är helt underbart " .
" Men jag valde att INTE belöna någon ( genom att köpa hans musik eller kläder eller stödja hans " konst " ) som jag tror omfamnar och sprider en ideologi som är skadlig för mitt samhälle .
Han är fri .
Det är vi med , tillade hon .
Innan showen meddelade rapparen på Twitter att han hade ändrat sitt namn och sa att han nu var " varelsen tidigare känd som Kanye West " .
Han är inte den första artisten att ändra sitt namn och följer i Diddys fotspår , även känd som Puff Daddy , Puffy och P Diddy .
Rapparkollegan , Snoop Dogg har kallat sig Snoop Lion och naturligtvis den avlidna musiklegenden Prince , ändrade sitt namn till en symbol och sedan till konstnären som tidigare var känd som Prince .
Dom för mordförsök efter knivskärning på restaurang i Belfast
En 45 @-@ årig man har anklagats för mordförsök efter att en man knivskars på en restaurang i östra Belfast på fredagen .
Händelsen inträffade i Ballyhackamore , sade polisen .
Svaranden förväntas infinna sig på Belfast Magistrates Court på måndagen .
Anklagelserna kommer att granskas av åklagarmyndigheten .
Game of Thrones @-@ stjärnan Kit Harington slår mot toxisk maskulinitet
Kit Harington är känd för sin svärdsvängande roll som Jon Snow i HBO:s våldsamma medeltida fantasy @-@ serie Game of Thrones .
Men skådespelaren , 31 , har uttalat sig negativt om stereotypen av machohjälten och säger att sådana roller på skärmen betyder att unga pojkar ofta känner att de måste vara tuffa för att respekteras .
I ett uttalande till Sunday Times Culture , sa Kit att han tror att " något har gått fel " och ifrågasatte hur man ska hantera problemet med toxisk maskulinitet under # MeToo @-@ eran .
Kit , som nyligen gifte sig med sin medskådespelare i Game of Thrones , Rose Leslie , även hon 31 , erkände att han känner " ganska starkt " för att ta itu med problemet .
" Jag känner personligen ganska starkt , just nu - var har vi gått fel med maskulinitet ? " , sa han .
" Hur har vi uppfostrat män med hänsyn till de problem vi ser nu ? "
Kit tror att TV delvis kan vara ansvarigt för ökningen av toxisk maskulinitet på grund av sina mycket maskulina karaktärer .
Han fortsatte " Vad är infött och vad är inlärt ?
Vad lärs ut på TV och på gatorna , som gör att unga pojkar känner att de måste vara på ett visst sätt för att vara man ?
Jag tror att det verkligen är en av de stora frågorna i vår tid - hur förändrar vi det ?
Det är tydligt att något har gått snett för unga män " .
I intervjun erkände han också att han inte skulle göra några Game of Thrones @-@ uppföljare när serien kommer till ett slut nästa sommar och säger att han är " klar med slagfält och hästar " .
Från november kommer Kit att spela i en nyinspelning av Sam Shepards True West som är berättelsen om en filmproducent och hans bror , som är en rånare .
Skådespelaren avslöjade nyligen att han tycker att mötet med sin fru Rose var den bästa erfarenheten från Game of Thrones .
" Jag träffade min fru tack vare serien , så på så sätt gav den mig min framtida familj och mitt framtida liv " , sa han .
Rose spelade Ygritte , som Kits karaktär Jon Snow förälskar sig i , i Emmys @-@ vinnande fantasy @-@ serien .
Paret gifte sig i juni 2018 på Leslies familjeägor i Skottland .
HIV / Aids : Kina rapporterar en 14 % ökning av nya fall
Kina har meddelat en ökning med 14 % av antalet medborgare som lever med hiv och aids .
Mer än 820 000 människor har drabbats i landet , säger hälsovårdsmyndigheterna .
Omkring 40 000 nya fall rapporterades bara under andra kvartalet 2018 .
De allra flesta nya fallen överfördes via sex och markerade en förändring från tidigare år .
Traditionellt sprids hiv snabbt genom vissa delar av Kina som ett resultat av infekterade blodtransfusioner .
Men antalet personer som smittas av HIV på detta sätt hade minskats till nästan noll , sade kinesiska hälsovårdsmyndigheter vid en konferens i Yunnanprovinsen .
Antalet personer som lever med hiv och aids i Kina har dock ökat med 100 000 personer från år till år .
HIV @-@ smitta genom samlag är en akut fråga i Kinas HBT @-@ community .
Homosexualitet avkriminaliserades i Kina år 1997 , men diskriminering av HBT @-@ personer sägs vara utbredd .
På grund av landets konservativa värderingar har studier uppskattat att 70 @-@ 90 % av männen som har sex med män förr eller senare kommer att gifta sig med kvinnor .
Många av smittofallen beror på otillräckligt skydd vid samlag i dessa relationer .
Kinas regering har sedan 2003 lovat universell tillgång till HIV @-@ medicin som en del av insatserna för att ta itu med problemet .
Maxine Waters nekar att personal läckt GOP @-@ senatorns uppgifter , skyler på " farliga lögner " och " konspirationsteorier "
Den amerikanska kongressledamoten Maxine Waters fördömde på lördagen påståenden om att en av hennes anställda hade lagt upp personuppgifter på tre republikanska amerikanska senatorer på deras Wikipedia @-@ sidor .
Los Angeles @-@ Demokraten hävdade att dessa påståenden spriddes av högerextremistiska webbplatser .
" Lögner , lögner och mer förkastliga lögner " , sade Waters i ett uttalande på Twitter .
Den släppta informationen innehöll enligt uppgift hemadresser och telefonnummer till senatorerna Lindsey Graham från South Carolina och Mike Lee och Orrin Hatch , båda från Utah .
Informationen uppkom online torsdag , upplagd av en okänd person på Capitol Hill under en senatpanels förhör om anklagelserna om sexuella övergrepp mot den nominerade kandidaten till Högsta domstolen , Brett Kavanaugh .
Läckan kom någon gång efter att de tre senatorerna ifrågasatte Kavanaugh .
Konservativa webbplatser som Gateway Pundit och RedState rapporterade att IP @-@ adressen som identifierar källan till inläggen var associerad med Waters kontor och släppte informationen om en medlem av Waters personal , rapporterade Hill .
" Detta ogrundade påstående är helt falskt och en absolut lögn " , fortsatte Waters .
" Min personal - vars identitet , personuppgifter och säkerhet har äventyras till följd av dessa bedrägliga och falska påståenden - var inte på något sätt ansvarig för läckan av denna information .
Detta ogrundade påstående är helt falsk och en absolut lögn " .
Waters uttalande fick snabbt kritik online , bland annat från Vita Husets tidigare press sekreterare Ari Fleischer .
" Detta förnekande är argt " , skrev Fleischer .
" Detta tyder på att hon inte har temperamentet att vara medlem av kongressen .
När någon anklagas för något de inte gjorde , får de inte vara arga .
De får inte vara trotsiga .
De får inte ifrågasätta ifrågasättarens motiv .
De måste vara lugna och sansade " .
Fleischer verkade försöka jämföra Waters reaktion med demokraternas kritik av domare Kavanaugh , som kritiker anklagade för att ha verkat vara arg under torsdagens förhör .
Omar Navarro , en republikansk kandidat som kandiderade för att avsätta Waters i mitten av mandatperioden uttryckte också sina tankar på Twitter .
" Stort om sant " , tweetade han .
I sitt uttalande sade Waters att hennes kontor hade varnat " lämpliga myndigheter och brottsbekämpande väsen för dessa bedrägliga krav .
" Vi kommer att se till att gärningsmännen kommer att avslöjas " , fortsatte hon " och att de kommer att hållas juridiskt ansvariga för alla sina handlingar som är destruktiva och farliga för alla mina anställda " .
Recension av Johnny English Strikes Again - kraftlös spionparodi av Rowan Atkinson
Det är nu tradition att leta efter Brexit @-@ betydelser i varje ny film med brittisk lutning , och detsamma verkar gälla för denna nyinspelning av den senaste Johnny English actionkomedin - en serie spionparodier som sparkades igång 2003 med Johnny English och fick nytt liv 2011 med Johnny English Reborn .
Kommer vass satir om hur uppenbart dåliga vi är att bli nationens nya exportvara ?
I alla fall har den den inkompetenta Johnny English med gummiansiktet fått sin licens att klanta till sake förnyats för andra gången - hans namn signalerar mer än något annat att han är en bred komisk skapelse avsedd för biopublik även i icke engelsktalande länder
Han är självklart den knäppa hemliga agenten , som trots sina bisarra anspråk på smoothieglamour har fått en liten bit av Clouseau , en gnutta Mr Bean och ett mått av killen från öppningsceremonin till OS i London 2012 .
Han är också ursprungligen baserad på den resenär och den internationella mystiska mannen som Atkinson en gång spelat i de nu glömda Barclaycard @-@ tv @-@ annonserna som skapar kaos vart han än går .
Det finns ett eller två fina ögonblick i den senaste JE @-@ filmen
Jag älskade när Johnny English närmar sig en helikopter klädd i en medeltida rustning och när rotorbladen en kort stund slog mot hans hjälm .
Atkinsons talang för fysisk komedi visas , men humorn känns ganska lågmäld och konstigt överflödig , speciellt eftersom de " seriösa " filmmärkena som 007 och Mission Impossible själva nu erbjuder komedi som en ingrediens .
Humorn känns som om den är anpassad för barn i stället för vuxna och för mig är Johnny English konstiga upptåg inte lika uppfinningsrika och fokuserade som Atkinsons stumfilmsbravader i rollen som Bean .
Det ständigt aktuella ämnet är nu att Storbritannien är i allvarliga problem .
En cyber @-@ hacker har infiltrerat Storbritanniens superhemliga webbnätverk av spioner , vilket avslöjar identiteterna av alla Storbritanniens agenter ute i fält , till agenten i tjänsts stora missnöje - en oerhört liten roll för Kevin Eldon .
Det blir det sista strået för en premiärminister som är en pompös och hårt ansatt figur , som redan lider av en fullständig kollaps av sin politiska popularitet : Emma Thompson gör sitt allra bästa med denna quasi @-@ Teresa @-@ May @-@ karaktär men manuset erbjuder inte mycket att jobba med .
Hennes underrättelserådgivare informerar henne om att när varje enskild aktiv spion är upptagen måste hon använda någon som gått i pension .
Och det betyder den stammande Johnny English i egen hög person , nu anställd som lärare i någon välbärgad institution , men som erbjuder inofficiella lektioner i konsten att arbeta undercover vid sidan av .
English skickades tillbaka till Whitehall för ett akut möte och återförenas med sin tidigare långlivade sidekick Bough , återigen spelad av av Ben Miller .
Bough är nu gift med en ubåtskapten , en jolly @-@ hockey @-@ sticks @-@ roll där Vicki Pepperdine är nära på bortkastad .
Så Batman och Robin är tillbaka efter det att allt gick så fruktansvärt fel på Her Majesty ' s Secret Service och stöter på Olga Kurylenkos vackra femme fatale Ophelia Bulletova .
Under tiden kommer premiärministern att falla hårt för den karismatiska techmiljardären , som hävdar att han kan lösa Storbritanniens datorbråk : den olyckliga Jason Volta , som spelas av Jake Lacy .
English och Bough börjar sin odyssé av farsartade upptåg : utklädda till servitörer , sätter de eld på en flashig fransk restaurang ; de skapar kaos när de smugglar sig ombord på Voltas lyxbåt ; och English utlöser ren anarki när han försöker använda ett VR @-@ headset för att bekanta sig med insidan av Voltas hus .
Det ligger säkerligen en hel del jobb bakom den sistnämnda sekvensen , men trots att filmen är både charmig och fartfylld , har den en air av barn @-@ TV kring sig .
Ganska måttligt allt som allt .
Och som med de andra Johnny English @-@ filmerna kan jag inte låta bli att tänka : Kan inte den brittiska filmindustrin ge Rowan Atkinson en roll som matchar hans talang ?
Labour förnekar att man utarbetar en plan för att britter ska arbeta en fyradagars vecka men få lön för fem dagar
Jeremy Corbyns parti Labour överväger en radikal plan som går ut på att britterna arbetar en fyra dagars vecka - men får betalt för fem .
Partiet vill enligt uppgift att företagsledare överlåter besparingar gjorda genom revolutionen i artificiell intelligens ( AI ) till arbetstagare genom att ge dem en extra ledig dag .
Det skulle se anställda njuta av en tre dagars helg - men behålla samma lön .
Enligt källor skulle idén " passa " med partiets ekonomiska agenda till förmån för arbetarna .
Att byta till en fyra dagars vecka har godkänts av fackorganisation Trades Union Congress som ett sätt för arbetstagare att dra fördel av ekonomiska förändringar .
En representant högre upp i Labor sa till The Sunday Times : En granskning av policyn förväntas offentliggöras före årets slut .
" Det kommer inte att ske på en dag , men en fyra dagars arbetsvecka är en strävan som passar in i partiets inställning till att balansera ekonomin till förmån för arbetaren samt partiets övergripande industriella strategi " .
Labour Party skulle inte vara den första som stöder en sådan idé , även partiet The Greens som lovade en fyra dagars arbetsvecka under sin valkampanj år 2017 .
Detta mål är dock inte påtecknad av Labour som helhet .
En talesman för Labour sade : " En fyradagars arbetsvecka är inte partiets policy och det är inget som partiet är överens om " .
Skuggkansler John McDonnell använde förra veckans Labour @-@ konferens för att kommunicera sin vision av en socialistisk revolution i ekonomin .
McDonnell sa att han var fast besluten att ta tillbaka makten från " ansiktslösa ledare " och " snyltare " på statliga företag .
Skuggkanslerens planer innebär också att de nuvarande aktieägarna i vattenföretag inte kan få tillbaka hela sin insats , eftersom en Labour @-@ regering kan göra " avdrag " på grund av vad de uppfattar har varit felaktiga handlingar .
Han bekräftade också planer på att sätta arbetstagare i företagsstyrelser och skapa så kallade Inclusive Ownership Funds där 10 procent av det privata företagets egna kapital lämnas över till dess anställda , som då står att få årliga utdelningar på upp till 500 pund .
Lindsey Graham och John Kennedy berättar i TV @-@ programmet " 60 minutes " om huruvida FBI:s utredning av Kavanaugh skulle kunna ändra deras åsikter
FBI:s utredning av anklagelser mot domare Brett Kavanaugh har försenat en slutlig omröstning om hans nominering till högsta domstolen med minst en vecka och lyfter frågan om huruvida byråns utredningar skulle kunna få några republikanska senatorer att ändra ställning i frågan .
I en intervju som sändes i söndags , frågade " 60 Minutes " korrespondent Scott Pelley de republikanska senatorerna John Kennedy och Lindsey Graham om huruvida FBI skulle kunna avslöja om någonting som skulle leda till att de ändrar åsikt .
Kennedy verkade mer öppen än sin kollega från South Carolina .
" Självklart " , sa Kennedy .
" Jag sa när jag gick in i utfrågningen , jag har pratat med domare Kavanaugh .
Jag ringde honom efter det att det hände , att påståendet kom ut , och sa : " Har du gjort det ? "
Han var bestämd , övertygad , otvetydig " .
Grahams röst verkar dock orubblig .
" Jag har redan bestämt mig angående Brett Kavanaugh och det skulle ta en dynamitanklagelse " , sa han .
" Dr . Ford , jag vet inte vad som hände , men jag vet det här : Brett förnekade det kraftigt " , tillade Graham , med hänvisning till Christine Blasey Ford .
" Och alla hon namnger kunde inte verifiera det .
Det var 36 år sen .
Jag ser inte att något nytt förändras " .
Vad är Global Citizen Festival och har det gjort något för att minska fattigdom ?
Denna lördag kommer New York att vara värd för Global Citizen Festival , en årlig musikhändelse som har en enormt imponerande uppställning av stjärnor som uppträder och ett lika imponerande uppdrag ; att bekämpa världsfattigdomen .
Nu under sitt sjunde år kommer Global Citizen Festival att se tiotusentals människor vallfärda till Central Parks Great Lawn , inte bara för att njuta av artister som Janet Jackson , Cardi B och Shawn Mendes , utan även för att öka medvetenheten om evenemangets verkliga mål : att bekämpa extrem fattigdom innan år 2030 .
Global Citizen Festival är , enligt ett uttalande från 2012 , en förlängning av Global Poverty Project , en internationell förespråksgrupp som hoppas kunna bekämpa fattigdom genom att öka antalet personer som aktivt kämpar mot den .
För att få en gratis biljett till evenemanget ( om du inte var redo att betala för en VIP @-@ biljett ) , skulle konsertgästerna utföra en serie uppgifter , eller " åtgärder " såsom volontärarbete , maila en världsledare , ringa eller på andra meningsfulla sätt bidra till att öka medvetenheten om målet att få slut på fattigdom .
Men hur framgångsrikt har Global Citizen varit med 12 år kvar för att nå sitt mål ?
Är idén att belöna människor med en gratis konsert ett genuint sätt att övertyga människor att agera , eller handlar det bara om så kallad " clicktivism " - människor som känner att de gör verklige skillnad genom att signera en online @-@ ansökan eller skriva ett tweet ?
Sedan 2011 uppger Global Citizen att man har registrerat mer än 19 miljoner " handlingar " från sina anhängare som kämpat för en mängd olika mål .
Det står att dessa åtgärder har bidragit till att sporra världsledare att tillkännage åtaganden och politik som motsvarar mer än 37 miljarder dollar , vilket kommer att påverka livet för mer än 2,25 miljarder människor år 2030 .
I början av 2018 citerade gruppen 390 åtaganden och tillkännagivanden som härrör från sina åtgärder , varav minst 10 miljarder dollar redan har betalats ut eller finansierats .
Gruppen uppskattar att de insamlade tillgångarna hittills har haft en direkt inverkan på nästan 649 miljoner människor över hela världen .
Några av de viktigaste åtagandena är The Power of Nutrition , ett partnerskap baserat i Storbritannien mellan investerare och aktörer som är engagerade i att " hjälpa barn att utvecklas till sin fulla potential " , lovande att ge Rwanda 35 miljoner dollar för att bidra till att bekämpa undernäring i området efter att ha fått mer än 4 700 tweets från globala medborgare .
" Med stöd från den brittiska regeringen , givare , nationella regeringar och globala medborgare , precis som du , kan vi göra sociala orättvisa som undernäring är till en fotnot i historien " , sade ambassadören för partnerskapet Tracey Ullman till folkmassan under en livekonsert i London i april 2018 .
Gruppen sade också att efter mer än 5000 åtgärder vidtagits som kräver att Storbritannien förbättrar kosten för mödrar och barn , tillkännagav regeringen finansiering av projektet , Power of Nutrition , som omfattar kostprogram som riktar sig till 5 miljoner kvinnor och barn .
Som svar på en av de vanliga frågorna på sin hemsida : " vad får dig att tro att vi kan bekämpa extrem fattigdom ? "
Svarade Global citizen : " Det kommer att bli en lång och svår väg - ibland kommer vi att falla och misslyckas .
Men , som de stora medborgerliga rättighets- och anti @-@ apartheidrörelserna innan oss , kommer vi att lyckas , för vi är starkare tillsammans .
Janet Jackson , the Weeknd , Shawn Mendes , Cardi B , Janelle Monáe är några av de artister som uppträder vid årets evenemang i New York , vars värdar är Deborra @-@ Lee Furness och Hugh Jackman .
USA skulle kunna använda sin flotta i en " blockad " för att hindra rysk energiexport anger inrikesministern
Regeringen kan " vid behov " tillgripa sin flotta för att förhindra ryska energiaktörer från att slå sig in på marknaderna , däribland i Mellanöstern , har amerikanska inrikesministern Ryan Zinke avslöjat , citerad av Washington Examinator .
Zinke påstod att Rysslands engagemang i Syrien - särskilt där det verkar på inbjudan från den legitima regeringen - är en förevändning för att utforska nya energimarknader .
" Jag tror att de är i Mellanöstern eftersom de vill sälja energi , precis som de gör i Östeuropa , Europas sydliga delar " , har han sagt .
Och enligt honom finns det sätt och medel att ta itu med det .
" USA har förmågan att , med vår flotta , se till att sjövägarna hålls öppna och , om nödvändigt , tillämpa blockad , för att se till att deras energi inte når marknaden " , sa han .
Zinke talade till deltagarna i evenemanget som anordnades av Consumer Energy Alliance , en ideell grupp som kallar sig för " energikonsumentens röst " i USA .
Han jämförde Washingtons tillvägagångssätt för att hantera Ryssland och Iran , och noterade att de verkligen är desamma .
" Det ekonomiska alternativet gentemot Iran och Ryssland är mer eller mindre att utnyttja och byta ut bränslen " , sade han , medan han hänvisade till Ryssland som en " dagsslända " med en ekonomi som är beroende av fossila bränslen .
Uttalanden kommer efter att Trump @-@ administrationen har haft som mål att öka exporten av sin flytande naturgas till Europa , för att ersätta Ryssland , det långt billigare alternativet för europeiska konsumenter .
I detta syfte försöker Trump @-@ administrationens tjänstemän , inklusive USA:s president Donald Trump , att övertyga Tyskland om att dra sig ur det " olämpliga " Nord Stream 2 @-@ pipelineprojektet , vilket enligt Trump gjorde Berlin till Moskvas " fånge " .
Moskva har upprepade gånger betonat att Nord Stream 2 @-@ rörledningen på 11 miljarder dollar , som ska dubbla den befintliga rörledningskapaciteten till 110 miljarder kubikmeter , är ett rent ekonomiskt projekt .
De hävdar att Washingtons motstånd mot projektet bara drivs av ekonomiska skäl och är ett exempel på illojal konkurrens .
" Jag tror att vi delar uppfattningen att energi inte kan vara ett verktyg för att utöva påtryckningar och att konsumenterna ska kunna välja leverantörerna " , sade Rysslands energiminister Alexander Novak efter ett möte med USA:s energisekreterare Rick Perry i Moskva i september .
Den amerikanska ståndpunkten fick bakslag från Tyskland , som har bekräftat sitt engagemang för projektet .
Tysklands ledande branschorganisation , Federation of German Industries ( BDI ) , har uppmanat USA att hålla sig borta från EU:s energipolitik och de bilaterala avtalen mellan Berlin och Moskva .
" Jag ogillar starkt att en tredje part stör vår energiförsörjning " , sade Dieter Kempf , chef för Federation of German Industries ( BDI ) efter ett möte mellan förbundskansler Angela Merkel och Rysslands president Vladimir Putin .
Elizabeth Warren kommer att ta en " ordentlig funderare " om hon ska ställa upp i presidentvalet 2020 , säger Massachusetts Senator
Massachusetts Senator Elizabeth Warren sade på lördag att hon skulle ta en " ordentlig funderare " kring hennes deltagande i presidentvalet efter USA:s mellanårsval .
Under ett rådhusmöte i Holyoke , Massachusetts , bekräftade Warren att hon skulle överväga att ställa upp som kandidat .
" Det är dags för kvinnor att ta sig till Washington och fixa vår trasiga regering och det inkluderar en kvinna på toppen " , sa hon enligt The Hill .
" Efter den 6 november kommer jag att ta en rejäl funderare på att kandidera till presidentposten " .
Warren vägde in på president Donald Trump under rådhusmötet och sa att han " tog detta land i fel riktning .
" Jag är djupt orolig över vad Donald Trump gör för vår demokrati " , sa hon .
Warren har varit frispråkig i sin kritik av Trump och hans kandidat till Högsta domstolen , Kavanaugh .
I en tweet på fredagen sade Warren " vi behöver naturligtvis en FBI @-@ utredning innan vi röstar " .
En omröstning som släpptes på torsdagen visade emellertid att en majoritet av Warrens egna anhängare inte trodde att hon skulle kandidera 2020 .
Femtioåtta procent av " troliga " Massachusettsväljare sade att senatorn inte borde kandidera , enligt en undersökning utförd av Suffolk University Political Research Center / Boston Globe .
Trettiotvå procent stödde kandidaturen .
Undersökningen visade mer stöd för en kandidatur av före detta guvernören Deval Patrick , med 38 procent för en potentiell kandidatur och 48 procent emot .
Andra högprofilerade demokratiska namn som diskuteras med avseende på en potentiell 2020 @-@ kandidatur inkluderar tidigare vicepresident Joe Biden och Vermonts Senator Bernie Sanders .
Biden sa att han skulle bestämma sig officiellt i januari , rapporterade Associated Press .
Sarah Palin citerar Track Palins PTSD vid Donald Trump rally
Track Palin , 26 , tillbringade ett år i Irak efter att ha tagit värvning i september .
Han greps och anklagades för våld i hemmet på måndagskvällen
" Vad min egen son går igenom , vad han går igenom nu när han är tillbaka , jag kan relatera till andra familjer som har erfarenhet av PTSD och en del av det trauma som våra soldater återvänder med " , sa hon till publiken vid ett samlingsmöte för Donald Trump i Tulsa , Oklahoma .
Palin kallade hans gripande för " elefanten i rummet " och sa om sin son och andra krigsveteraner att " de kommer tillbaka som andra människor , de kommer tillbaka härdade , de kommer tillbaka och undrar om det finns respekt för det som deras kollegor , soldater och flygare och alla andra medlemmar i militären , har gett landet . "
Han greps på måndagen i Wasilla , Alaska och anklagades för våld i hemmet gentemot en kvinna , försök till hindrande av en rapport om våld i hemmet och vapeninnehav i berusat tillstånd , enligt Dan Bennett , en talesman för Wasilla Police Department .
18 stater , samt District of Columbia stöder ifrågasättandet av en ny asylpolitik
Arton stater och District of Columbia stöder en rättslig prövning riktad mot en ny amerikansk politik som förnekar asyl till offer som flyr gängrelaterat våld eller våld i hemmet .
Företrädare från de 18 staterna och distriktet inlämnade en friend @-@ of @-@ the @-@ court @-@ ansökan på fredagen ​ ​ i Washington för att stödja en asylsökande som utmanar policyn , rapporterade NBC News .
Fullständigt namn på käranden i ärendet Grace v . Sessions som American Civil Liberties Union inlämnade i augusti mot policyn har inte avslöjats .
Hon sa att hennes partner " och hans våldsamma gängmedlemsöner " , misshandlade henne , men amerikanska tjänstemän nekade hennes asylansökan den 20 juli .
Hon fängslades i Texas .
Staternas advokater som stöder Grace beskrev El Salvador , Honduras och Guatemala , länder som producerar ett stort antal asylsökande , som nationer som står inför stora problem med gäng och våld i hemmet .
Den nya amerikanska asylpolitiken ändrade ett beslut av immigrationsmyndigheterna från 2014 som gjorde det möjligt för olagliga invandrare att söka asyl för att fly från våld i hemmet .
District of Columbia Attorney General Karl Racine sade i ett uttalande på fredagen ​ ​ att den nya politiken " ignorerar decennier av statlig , federal och internationell rätt " .
" Federal lag kräver att alla asylansökningar ska bedömas baserat på särskilda fakta och omständigheter som fordran gäller , och en sådan bestämmelse strider mot den principen " , enligt friend @-@ of @-@ the court @-@ rapporten .
Advokater hävdade vidare i rapporten att politiken som förnekar invandrarnas inträde skadar den amerikanska ekonomin , och argumenterar att de är mer benägna att bli entreprenörer och " leverera nödvändig arbetskraft " .
Justitieministern Jeff Sessions beordrade i juni domare i asylfall att inte längre bevilja asyl till offer som flydde våld i hemmet och gängvåld .
" Asyl är tillgängligt för dem som lämnar sitt hemland på grund av förföljelse eller rädsla på grund av ras , religion , nationalitet eller medlemskap i en viss social grupp eller politisk åsikt " sa Sessions när policyn tillkännagavs 11 juni .
Asyl var aldrig menat att lindra alla problem - även alla allvarliga problem - som människor står inför varje dag över hela världen .
Desperata räddningsinsatser i Palu när dödssiffran fördubblas i jakten på överlevande
För de överlevande såg situationen allt dystrare ut .
" Det känns väldigt spänt " , sade den 35 @-@ årige mamman Risa Kusuma , som tröstade sin febriga pojke i ett evakueringscenter i staden Palu .
" Ambulansen hämtar döda kroppar hela tiden .
Rent vatten är en bristvara " .
Invånarna sågs återvända till sina förstörda hem , rotandes genom vattenskadade ägodelar och försökte rädda allt de kunde hitta .
Hundratals människor skadades och sjukhus , som skadats i jordbävningen på 7.5 var överfulla .
Några av de skadade , inklusive Dwi Haris , som drabbades av en bruten rygg och axel , vilade utanför sjukhuset Palu ' s Army Hospital , där patienterna behandlades utomhus på grund av fortsatt starka efterskalv .
Med tårfyllda ögon berättade han att den våldsamma jordbävningen skakade rummet på hotellets femte våning som han delade med sin fru och dotter .
" Vi hann inte fly .
Jag pressades in i murens ruiner , tror jag " , berättade Haris för Associated Press och tillade att hans familj var i stan för ett bröllop .
" Jag hörde min fru skrika på hjälp , sen blev det tyst .
Jag vet inte vad som hände med henne och mitt barn .
Jag hoppas att de är i säkerhet " .
USA:s ambassadör anklagar Kina för " mobbning " med " propagandaannonser "
En vecka efter att en officiell kinesisk tidning publicerade en fyrsidig annons i en amerikansk dagstidning om de ömsesidiga fördelarna av handeln mellan USA och Kina , anklagade den amerikanska ambassadören till Kina att Peking använde den amerikanska pressen för att sprida propaganda .
USA:s President Donald Trump hänvisade förra onsdagen till att China Daily betalade ett tillskott i Des Moines Register - staten Iowas bäst säljande tidning - efter att ha anklagat Kina för att försöka medverka i USA:s 6:e kongressval , något som Kina förnekar .
Trumps anklagelse att Peking försökte blanda sig i amerikanska val markerade vad amerikanska tjänstemän berättade för Reuters var är en ny fas i en eskalerande kampanj från Washington ämnad att sätta press på Kina .
Även om det är normalt för utländska regeringar att använda reklam för att främja handel , är Peking och Washington för tillfället låsta i ett eskalerande handelskrig med höjda tariffer på varandras importer .
Kinas vedergällningstariffer tidigt i handelskriget utformades för att drabba exportörer i stater som Iowa som stöder Trumps republikanska parti , detta enligt kinesiska och amerikanska experter .
Terry Branstad , USA:s ambassadör i Kina och den tidigare långvariga guvernören i Iowa , en stor exportör av jordbruksprodukter till Kina , sa att Peking hade skadat amerikanska arbetare , bönder och företag .
Kina , skrev Branstad i en debattartikel i söndagens Des Moines Register , " fördubblar nu mobbningen genom att lägga ut propagandaannonser i vår egen fria press " .
" Kinas regering använder sig av Amerikas kära tradition av yttrandefrihet och en fri press för att sprida propagandan till genom att publicera betalda reklamannonser i Des Moines Register " , skrev Branstad .
" I kontrast , i tidningskiosken på gatan här i Peking hittar du ett begränsat antal avvikande röster och kommer inte att se någon sann avspegling av de olika åsikter som det kinesiska folket kan ha om Kinas oroliga ekonomi , eftersom media styrs med järnhand av det kinesiska kommunistpartiet , " skrev han .
Han tillade att " en av Kinas mest framstående tidningar nobbade erbjudandet att publicera " hans artikel , även om han inte sa vilken tidning .
Republikaner skrämmer bort kvinnliga väljare inför mellanårsvalet genom Kavanaugh @-@ fiaskot , varnar analytiker
Eftersom många topprepublikaner försvarar högsta domstolens nominerade Brett Kavanaugh som står inför flera anklagelser om sexuella övergrepp , har analytiker varnat för att det kommer ske ett bakslag , särskilt från kvinnor , under det kommande valet .
Känslorna kring detta har varit extremt höga , och de flesta republikaner har redan visat var de står i valet .
Det går inte att vrida tillbaka klockan , säger Grant Reeher , professor i statsvetenskap vid Syracuse Universitys Maxwell School , till The Hill i en artikel som publicerades i lördags .
Reeher sa att han tvivlar på senator Jeff Flakes ( R @-@ Arizona ) sista försök till en en FBI @-@ utredning kommer att räcka för att lugna arga väljare .
" Kvinnor kommer inte att glömma vad som hände igår - de kommer inte att glömma det imorgon och inte i november " , säger Karine Jean @-@ Pierre , en seniorrådgivare och nationell taleskvinna för den progressiva gruppen MoveOn på fredagen , enligt tidningen Washington , DC .
På fredag ​ ​ morgon skanderade de demonstrerande " November kommer ! " när de demonstrerade i hallen till senatbyggnaden när republikanerna som kontrollerar domstolskommittén valde att gå vidare med Kavanaughs nominering trots vittnesmålet från Dr . Christine Blasey Ford , rapporterade Mic .
" Demokratisk entusiasm och motivation kommer att gå i taket " , berättade Stu Rothenberg , en neutral politisk analytiker , för nyhetssajten .
" Folk säger att det redan varit högt , det är sant .
Men det kunde vara högre , särskilt bland ännu obestämda kvinnliga väljare i förorterna och yngre väljare , 18- till 29 @-@ åringar , som , trots att de inte gillar presidenten , ofta inte röstar " .
Redan innan Fords offentliga vittnesmål med anklagelser om sexuella övergrepp mot den nominerade kandidaten till högsta domstolen , föreslog analytiker att ett bakslag kunde följa om republikanerna pressade igenom bekräftelsen .
" Det här har blivit en förvirrad röra för GOP " , sade Michael Steele , tidigare ordförande för den republikanska nationella kommittén , i början av förra veckan , enligt NBC News .
" Det handlar inte bara om kommitténs omröstning eller slutomröstningen eller om Kavanaugh kommer igenom , det handlar också om hur republikaner har hanterat detta och hur de har behandlat henne " , påpekade Guy Cecil , chef för Priorities USA , en grupp som hjälper demokratiska valkampanjer , för nyhetskanalen .
Men amerikanerna i allmänhet verkar vara delade över vem de ska tro på i kölvattnet av Fords och Kavanaughs vittnesmål , och den senare verkar vara den de tror mest på .
En ny opinionsundersökning från YouGov visar att 41 procent av respondenterna definitivt eller troligen trodde på Fords vittnesbörd , medan 35 procent sa att de definitivt eller troligen trodde på Kavanaugh .
Dessutom sa 38 procent att de tyckte att Kavanaugh troligen eller definitivt ljugit under sitt vittnesbörd , medan bara 30 procent sa detsamma om Ford .
Efter påtryckningar från Flake , undersöker FBI för närvarande de påståenden som Ford har framfört , liksom de från minst en annan anklagare , Deborah Ramirez , rapporterade The Guardian .
Ford vittnade inför senatens domstolskommitté under ed i förra veckan att Kavanaugh våldsamt angrep henne vid 17 års ålder .
Ramirez hävdar att den kandidaten till högsta domstolen exponerade sina könsorgan för henne medan de deltog i en fest under deras tid som studenter vid Yale på 1980 @-@ talet .
Uppfinnaren av World Wide Web planerar att starta ett nytt internet för att konkurrera med Google och Facebook
Tim Berners @-@ Lee , uppfinnaren av World Wide Web , lanserar en startup som syftar till att konkurrera med Facebook , Amazon och Google .
Teknologilegendens senaste projekt , Inrupt , är ett företag som bygger sig på Berners @-@ Lees open source @-@ plattform Solid .
Solid tillåter användare att välja var deras data lagras och vilka personer som får tillgång till vilken information .
I en exklusiv intervju med Fast Company skämtade Berners @-@ Lee att avsikten bakom Inrupt är " världsdominans " .
" Vi måste göra det nu " , sa han om startup @-@ företaget .
" Det är ett historiskt ögonblick " .
Appen använder Solids teknik för att tillåta människor att skapa sin egen " personal online data store " eller en POD .
Den kan innehålla kontaktlistor , att göra @-@ listor , kalender , musikbibliotek och andra personliga och professionella verktyg .
Det är som om Google Drive , Microsoft Outlook , Slack och Spotify alla är tillgängliga i en webbläsare samtidigt .
Det som är unikt med den personliga online @-@ datalagringen är att det är helt upp till användaren vem som kan få tillgång till vilken typ av information .
Företaget kallar det " personligt bemyndigande genom data " .
Idén med Inrupt , enligt företagets VD John Bruce , är att företaget ska ta med resurser , processer och lämpliga färdigheter för att göra Solid tillgängligt för alla .
Företaget består för närvarande av Berners @-@ Lee , Bruce , en säkerhetsplattform som köptes av IBM , en del programutvecklare som ska arbeta med projektet och en grupp volontärkodare .
Från och med denna vecka kan teknikutvecklare runt om i världen skapa egna decentraliserade appar med hjälp av de verktyg som finns tillgängliga på Inrupt @-@ webbplatsen .
Berners @-@ Lee sa att han och hans team inte pratar med " Facebook och Google om huruvida man ska introducera en komplett förändring där alla affärsmodeller ställs på högkant över en natt .
" Vi ber dem inte om tillåtelse " .
I ett inlägg på Medium som publicerades på lördagen , skrev Berners @-@ Lee att Inrupts uppdrag är att tillhandahålla kommersiell energi och ett ekosystem för att skydda integriteten och kvaliteten på den nya webben som skapas av Solid .
1994 omvandlade Berners @-@ Lee Internet när han etablerade World Wide Web Consortium vid Massachusetts Institute of Technology .
Berners @-@ Lee har de senaste månaderna varit en inflytelserik röst i debatten om nätneutralitet .
Även under lanseringen av Inrupt kommer Berners @-@ Lee att fortsätta vara grundare och chef för World Wide Web Consortium , Web Foundation och Open Data Institute .
" Jag är mycket optimistisk inför den här nya eran på webben " , tillade Berners @-@ Lee .
Bernard Vann : Präst belönad med Viktoria @-@ kors under första världskriget firas
Den enda prästen inom engelska kyrkan som belönades med ett Victoria @-@ kors under första världskriget firas nu i sin hemstad 100 år senare .
Lt Col Reverend Bernard Vann fick utmärkelsen för sitt agerande under attacken på Bellenglise och Lehaucourt den 29 september 1918 .
Han dödades dock av en prickskytt fyra dagar senare och fick aldrig veta att han hade tilldelats den brittiska militärens mest prestigefyllda pris .
En minnessten avtäcktes av hans två barnbarn under en parad i Rushden , Northamptonshire , på lördagen .
Ett av hans barnbarn , Michael Vann , sa att det var " briljant symboliskt " , att stenen skulle avslöjas exakt 100 år efter det att hans farfar belönats med priset .
Enligt London Gazette ledde Lt Col Vann den 29 september 1918 sin bataljon över Canal de Saint @-@ Quentin " genom en mycket tjock dimma och under tung eld från fält- och maskingevär " .
Han rusade senare upp till skottlinjen och ledde med " stor tapperhet " linjen framåt innan han ensam avgjorde striden .
Lt Col Vann dödades av en tysk prickskytt den 4 oktober 1918 - lite mer än en månad innan krigets slut .
Michael Vann , 72 , sa att hans farfars handlingar var " något som jag vet att jag aldrig kunde leva upp till , men något jag är mycket ödmjuk inför " .
Han och hans bror Dr James Vann lade också ner en krans efter paraden , som leddes av Brentwood Imperial Youth Band .
Michael Vann sa att han " kände sig mycket hedrad att spela en roll i paraden " och tillade att " en äkta hjältes mod demonstreras av det stöd som kommer att ges av många människor " .
MMA fans stannade uppe hela natten för att titta på Bellator 206 och fick istället se Greta Gris
Föreställ dig det här , du har stannat upp hela natten för att se Bellator 206 bara för att bli nekad att titta på huvudevenemanget .
Showen från San Jose innehöll 13 matcher , inklusive sex på huvudkortet och visades live på natten i Storbritannien på kanal 5 .
Klockan 06 : 00 , precis som Gegard Mousasi och Rory MacDonald förberedde sig för att möta varandra , överraskades de brittiska tittarna när programmet plötsligt ändrades till Greta Gris .
Många var föga imponerade efter att de hade hållit sig vakna till de tidiga morgontimmarna för att titta på matchen .
En fan på Twitter beskrev programändringen till ett tecknat barnprogram som " ett sjukt skämt " .
" Det var regeringens beslut att innehållet inte var lämpligt så tidigt på morgonen , så de var tvungna att byta till barnprogram " , sa Dave Schwartz , Bellators vice vd för marknadsföring och kommunikation när han frågades om sändningen .
" Greta gris , ja "
Bellators VD Scott Coker sa att de kommer att arbeta med sin schemaläggning för att bättre inkludera brittiska tittare i framtiden .
" Jag tror att vi kommer att kunna hitta en lösning vad gäller reprisen , sa Coker .
" Men det är sex på morgonen på en söndag där och vi kommer inte kunna lösa det här till söndag vår tid , måndag deras tid .
Men vi jobbar på det .
Tro mig , programbytet upprörde många .
Vi försökte åtgärda det , vi trodde att det rörde sig om ett tekniskt fel .
Men det var i själva verket en statlig fråga .
Jag kan lova att det inte kommer att hända nästa gång .
Vi kommer att visa fem matcher i stället för sex - som vi normalt gör . Vi tog oss vatten över huvudet i vår strävan efter att tillfredsställa fansen .
Det är en olycklig situation " .
Desert Island Discs : Tom Daley kändes " underlägsen " på grund av sexualitet
Den olympiska dykaren Tom Daley säger att kände sig underlägsen sina kamrater under sin uppväxt på grund av sin sexualitet - men det sporrade honom också till att bli framgångsrik .
24 @-@ åringen sa att han inte insåg att han inte var som alla andra förrän han gick på gymnasiet " .
När han talade i den första Radio 4 Desert Island Discs presenterad av Lauren Laverne sa han att han talade om homosexuellas rättigheter för att ge andra " hopp " .
Han sa också att han brydde sig mindre om att vinna OS efter att blivit förälder .
Den populära showens ordinarie programledaren , Kirsty Young , har tagit ledigt några månader på grund av sjukdom .
Under sitt engångsuppträdande på Lavernes första program berättar Daley hur han han kände sig " mindre värd " än andra under sin uppväxt , för att " det inte var inte socialt acceptabelt att tycka om pojkar och tjejer " .
Han sa : " Den här känslan av att känna mig mindre värd och känna mig annorlunda har varit en verklig källa till kraften och styrkan att lyckas " .
Han ville bevisa att han var " någon " , sa han , så att han inte svek alla när de så småningom fick reda på hans sexualitet .
Den tvåfaldige olympiske bronsmedaljören har blivit en högprofilerad förespråkare för HBT @-@ rättigheter och utnyttjade sitt framträdande vid årets Commonwealth Games i Australien för att övertyga fler länder att avkriminalisera homosexualitet .
Han sa att han tog till orda eftersom han kände sig ha haft turen att kunna leva öppet utan begränsningar och ville ge andra " hopp " .
Den trefaldige världsmästaren sa att hans förälskelse i en man - den amerikanska filmmakaren Dustin Lance Black , som han träffade 2013 - " kom som en överraskning " .
Daley gifte sig med den 20 år äldre Oscarsvinnaren förra året men han sa att åldersskillnaden aldrig hade varit ett problem .
" När du går igenom så mycket i en sådan ung ålder " - han deltog i sitt första OS som 14 @-@ åring och hans far dog av cancer tre år senare - sa han att det var svårt att hitta någon i samma ålder med liknande livserfarenhet .
Paret blev föräldrar i juni till en son vid namn Robert Ray Black @-@ Daley , och Daley sa att hans " hela livsperspektiv " hade förändrats .
" Om du hade frågat mig förra året handlade det bara om att vinna guld , sa han .
" Men vet du , det finns större saker än olympiska guldmedaljer .
Min guldmedalj är Robbie " .
Hans son bär samma namn som hans far Robert , som dog 2011 vid 40 års ålder efter att ha diagnostiserats med hjärncancer .
Daley sa att pappa inte accepterade att han skulle dö och en av de sista sakerna som han hade frågat om var om de fått sina biljetter till olympiska spelen i London 2012 - där han ville sitta på första raden .
" Jag kunde inte säga till honom : du kommer inte att kunna sitta på främre raden pappa " sa han .
" Jag höll hans hand när han slutade andas och det var inte förrän han faktiskt hade slutat andas och han var död som jag slutligen erkände att han inte var oövervinnerlig " , sa han .
Året därpå tävlade Daley vid OS 2012 och vann brons .
" Jag visste bara att det här var det jag hade drömt om hela mitt liv - att dyka framför en hemmapublik på en olympisk arena , det fanns ingen bättre känsla " , sa han .
Det inspirerade också hans första låtval - Proud av Heather Small - en låt som hade följt honom fram till OS och som fortfarande gav honom rysningar .
Desert Island Discs sänds på BBC Radio 4 på söndag kl. 11 : 15 BST .
Mickelson ur form på bänken under lördagens Ryder Cup
Amerikanen Phil Mickelson kommer slå rekord på söndag när han spelar sin 47:e Ryder Cup @-@ match , men då måste han fixa formen för att undvika en olycklig milstolpe .
Mickelson , som spelade för 12:e gången i rad , bänkades av kapten Jim Furyk för lördagens fourballs och foursomes .
I stället för att vara i händelsernas centrum , som han ofta har varit för USA , tillbringade den femfaldige vinnaren sin dag mellan att agera hejaklack och att träna på sitt spel i hopp om att få en chans att visa upp sin förmåga .
Han har aldrig varit den rakaste av drivers , inte ens på toppen av sin karriär och 48 @-@ åringen är inte i form inför den tuffa banan på Le Golf National , där den långa ruffen ofta straffar missar hårt .
Det är inte bara banan som avskräcker , i den nionde matchen på söndag möter Mickelson mästaren Francesco Molinari , som tillsammans med novisen Tommy Fleetwood vunnit alla fyra matcherna denna vecka .
Om amerikanerna , som ligger 4 poäng under inför de 12 singelmatcherna har medvind i starten , kan Mickelsons match vara helt avgörande .
Furyk uttryckte förtroende för sin spelare , inte för att han kunde säga mycket annat .
" Han förstod helt den roll som han hade idag , gav mig en klapp på ryggen och lade armen om mig och sa att han skulle vara redo imorgon " , sa Furyk .
" Hans självförtroende är det inget fel på .
Han är en kändis och han har tillfört så mycket till dessa lag under tidigare säsonger och under den gångna veckan .
Jag trodde förmodligen inte att han skulle klara av att spela två matcher .
Jag trodde han skulle klara mer , men nu är det som det är och vi får nöja oss med det .
Han vill vara där ute , precis som alla andra "
På söndagen passerar Mickelson Nick Faldo ' s rekord för flest Ryder Cup @-@ matcher spelade .
Det kan markera slutet på en Ryder Cup @-@ karriär som aldrig helt levt upp till höjderna i hans individuella resultat .
Mickelson har 18 segrar , 20 förluster och sju halvor , men Furyk sa att hans närvaro medfört andra kvaliteter laget .
" Han är rolig , han är sarkastisk , kvick , gillar att skämta med människor och han är en bra kille att ha i laget " , förklarade han .
" Jag tror också att de yngre spelarna tyckte det var roligt att spela mot honom den här veckan , vilket var kul att se .
Han tillför så mycket mer än bara spel " .
Europakaptenen Thomas Bjorn vet att den stora ledningen snart kan vara ett minne blott
Thomas Bjorn , den europeiska kaptenen , vet av erfarenhet att en betydande ledning i sista dagens singlar i Ryder Cup snabbt kan förändras till en obehaglig upplevelse .
Dane gjorde sin debut i 1997 års match på Valderrama , där ett lag under Seve Ballesteros ledning höll en fem @-@ poängs fördel över amerikanerna men som slutligen vann med minsta möjliga marginal med resultatet 14 ½ - 13 ½ .
" Man påminner dig om att vi ledde stort på Valderrama , vi ledde stort på Brookline där vi förlorade , och i Valderrama , där vi vann med nöd och näppe " , sa Bjorn ( på fotot ) efter att ha sett 2018 års klass vinna 5 @-@ 3 både i fredags ​ ​ och igår och leder med 10 @-@ 6 på Le Golf National .
Så historien kommer att bevisa för mig och alla i laget att detta inte är över .
Imorgon ger vi allt .
Går ut och gör allt rätt .
Detta är inte över förrän vi ser poängen på tavlan .
Vår målsättning är att försöka vinna denna pokal och det är där vårt fokus ligger .
Jag har sagt det hela tiden , jag fokuserar på de 12 spelare som finns på vår sida , men vi är väl medvetna om vad som väntar på andra sidan - de bästa spelarna i världen " .
Björn var nöjd med sina spelares prestationer på en tuff golfbana och tillade : " Jag skulle aldrig klara av detta själv .
Imorgon väntar nya utmaningar .
I morgon är det de enskilda prestationerna som gäller och det är en helt annan sak .
Det är kul att vara ute med en partner när det går bra , men när du är därute på egen hand , så testas din kapacitet som golfspelare fullt ut .
Det är budskapet som du behöver förmedla till spelarna , att få ut det bästa av sig själv imorgon .
Nu lämnar du din partner bakom dig och han måste också gå och få ut det bästa av sig själv " .
I motsats till Björn , kommer motståndaren Jim Furyk vilja att spelarna presterar bättre individuellt än de gjorde som partners , undantaget Jordan Spieth och Justin Thomas , som kammade hem tre poäng av fyra .
Furyk själv har varit på båda sidor av stora omvändningar under sista dagarna i en tävling , både i det vinnande laget i Brookline innan han slutade som förlorare när Europa körde " Miracle at Medinah " .
" Jag kommer ihåg vartenda jävla ord av det " , sa han som svar när han blev tillfrågad hur Ben Crenshaw , kaptenen 1999 , hade samlat sina spelare inför den sista dagen .
" Vi har 12 viktiga matcher imorgon , men man skulle vilja gå ut lika snabbt som på Brookline , som på Medinah .
När tempot kommer igång åt ena hållet blir det mycket press på dessa mellanmatcher .
Vi gjorde vår uppställning och placerade killarna som vi ville för att , du vet , skapa lite magi imorgon " .
Thomas fick uppgiften att försöka leda kampen och möter Rory McIlroy i toppmatchen , medan Paul Casey , Justin Rose , Jon Rahm , Tommy Fleetwood och Ian Poulter möter de andra européerna i översta halvan av ordningen .
" Jag gick med den här gruppen av killar i den här ordningen eftersom jag tycker att den räcker hela vägen " , sa Bjorn om sina singelval .
Tysklands nya krigsskepp senareläggs igen
Den tyska flottans nyaste fregatt skulle ha sjösatts 2014 för att ersätta krigsfartyg från det kalla krigets tid , men det kommer inte att sjösättas förrän åtminstone nästa år på grund av felaktiga system och höga kostnader , rapporterade lokala medier .
Idriftsättning av " Rheinland @-@ Pfalz " , ledskeppet för de helt nya Baden @-@ Wuerttemberg @-@ fregatterna , har nu skjutits upp till första halvåret 2019 , enligt Die Zeit @-@ tidningen som citerar en militär talesman .
Fartyget borde ha anslutit sig till flottan redan 2014 , men de problem som uppstod efter leveransen var ödesdigert för det ambitiösa projektet .
De fyra fartygen i Baden @-@ Wuerttemberg @-@ klass som flottan beställde 2007 kommer att ersätta de åldrande Bremen @-@ fregatterna .
De kommer att innehålla en kraftfull kanon , en rad luftvärns- och sjömålsmissiler , liksom vissa smygtekniker , såsom reducerad radar , infraröd och akustisk signatur .
Andra viktiga funktioner inkluderar längre underhållsperioder - det borde vara möjligt att stationera de nyaste fregatterna i upp till två år utan kontakt med hemmahamnar .
Men kontinuerliga förseningar innebär att de banbrytande krigsfartygen - som tillåter Tyskland att projektera makt utomlands - redan är föråldrade när de tas i drift , skriver Die Zeit .
Den ödesdigra F125 @-@ fregatten skapade rubriker förra året , då den tyska flottan officiellt vägrade att sätta fartyget i drift och returnerade det till Blohm & Voss varv i Hamburg .
Detta var första gången som flottan returnerat ett skepp till en skeppsbyggare efter leverans .
Lite var känt om orsakerna till returen , men tyska medier angav ett antal viktiga " mjukvaru- och maskinvarufel " som gjorde krigsskeppet värdelöst om det användes på ett stridsuppdrag .
Brister i programvaran var särskilt viktiga eftersom fartyg i Baden @-@ Wuerttemberg @-@ klassen kommer att drivas av en bemanning på cirka 120 sjömän - bara hälften av besättningen på äldre fregatter i Bremen @-@ klassen .
Det framkom också att fartyget har en betydande övervikt , vilket leder till försämrad prestanda och begränsar marinens förmåga att utföra framtida uppgraderingar .
Den 7 000 ton tunga " Rheinland @-@ Pfalz " antas vara dubbelt så tungt som likartade fartyg som användes av tyskarna under andra världskriget .
Bortsett från felaktig hårdvara , blir också hela projektets prislapp - inklusive utbildning av besättningen - ett problem .
Den sägs ha uppgått till svindlande 3,1 miljarder euro ( 3,6 miljarder dollar ) - jämfört med 2,2 miljarder euro i startskedet .
Problem som drabbar de nyaste fregatterna blir särskilt viktiga i ljuset av de senaste varningarna om att Tysklands sjömakt minskar .
Tidigare i år erkände Hans @-@ Peter Bartels , chef för det tyska parlamentets försvarskommitté , att flottan faktiskt " börjar få brist fullt utrustade fartyg " .
Tjänstemannen sade att det rör sig om ett växande problem , eftersom gamla fartyg avvecklas men inga ersättningsfartyg tillhandahölls .
Han beklagade att ingen av fregatterna i Baden @-@ Wuerttemberg @-@ klassen kunde ansluta sig till marinen .
National Trust tjuvlyssnar till fladdermössens hemliga liv
Ny forskning som utförs på en fastighet i de skotska högländerna syftar till att avslöja hur fladdermöss använder landskapet i sin jakt på mat .
Vi hoppas att resultaten kommer att kasta nytt ljus över beteendet hos unika flygande däggdjur och bidra till att styra framtida bevarandeaktiviteter .
Studien , utförd av forskare vid National Trust for Scotland , kommer att följa syd- och dvärgpipistrell samt bruna långörade och Daubenton fladdermöss på Inverewe Gardens i Wester Ross .
Särskilda inspelare kommer att placeras på viktiga platser runt fastigheten för att spåra fladdermusaktiviteter under hela säsongen .
NHS @-@ personal och volontärer kommer också att genomföra mobila undersökningar med hjälp av handhållna detektorer .
Expertljudanalys av alla inspelningar kommer att fastställa frekvensen av fladdermusljud och vilka arter som gör vad .
En livsmiljökarta och rapport kommer då att produceras för att skapa en detaljerad områdesbild av deras beteende .
Rob Dewar , naturvårdsrådgivare för NTS , hoppas att resultaten kommer att avslöja vilka områden av livsmiljö som är viktigast för fladdermössen och hur de används av var och en av arterna .
Denna information kommer att bidra till att bestämma fördelarna med livsmiljöhanteringsarbete såsom skapande av ängar och hur man bäst kan upprätthålla skogsmarker för fladdermöss och andra relaterade arter .
Fladdermuspopulationer i Skottland och i Storbritannien har minskat avsevärt under det senaste århundradet .
De hotas av byggnads- och utvecklingsarbete som påverkar bon och förlust av livsmiljöer .
Vindturbiner och belysning kan också utgöra en risk , liksom flygplan och vissa kemiska behandlingar av byggmaterial samt attacker från huskatter .
Fladdermöss är faktiskt inte blinda .
Men på grund av deras nattliga jaktvanor är deras öron mer användbara än deras ögon när det gäller att fånga byten .
De använder en sofistikerad eko @-@ lokaliseringsteknik för att hitta insekter och hinder i sin flygväg .
NTS , som ansvarar för vården av mer än 270 historiska byggnader , 38 viktiga trädgårdar och 76.000 hektar mark runt om i landet , tar fladdermöss på stort allvar .
Organisationen har tio utbildade experter , som regelbundet utför undersökningar , granskar bon och ibland utför räddningsoperationer .
Organisationen har även etablerat Skottlands första och enda dedikerade fladdermusreserv på Threave Estate i Dumfries och Galloway , hem för åtta av Skottlands tio fladdermusarter .
Egendomsförvaltaren David Thompson säger att egendomen är det idealiska området för dem .
" Här på Threave har vi ett bra område för fladdermöss " , sa han .
" Vi har de gamla byggnaderna , massor av veteranträd och en mängd gynnsamma livsmiljöer .
Men det finns mycket om fladdermöss som fortfarande är okänt , så det arbete vi gör här och på andra egendomar hjälper oss att förstå mer om vad de behöver för att trivas .
Han betonar vikten av att söka efter fladdermöss innan man utför underhåll inom fastigheter , eftersom det är möjligt att oavsiktlig förstörelse av ett enda bo skulle kunna döda upp till 400 honor och unga , och eventuellt utplåna en hel population .
Fladdermöss är fridlysta och det är olagligt att döda , besvära eller störa dem eller förstöra deras bon .
Elisabeth Ferrell , skotsk officer för Bat Conservation Trust , har uppmuntrat allmänheten att hjälpa till .
Hon sa : " Vi har fortfarande mycket att lära oss om våra fladdermöss och för många av våra arter vet vi inte hur deras populationer mår " .
Ronaldo avvisar våldtäktsdom medans hans advokater hotar att stämma den tyska tidningen
Cristiano Ronaldo har kallat våldtäktsanklagelserna mot honom för " falska nyheter " och säger att folk " vill marknadsföra sig " genom att använda hans namn .
Hans advokater kommer att stämma den tyska tidningen Der Spiegel , som publicerade påståendena .
Portugals och Juventus forward har anklagats för att ha våldtagit en amerikansk kvinna , Kathryn Mayorga , på ett hotell i Las Vegas 2009 .
Han påstås ha betalat henne 375,000 $ för att hålla tyst om händelsen , rapporterade Der Spiegel på fredagen .
I en Live @-@ video på Instagram slog Ronaldo ( 33 ) ifrån sig rapporterna som " falska nyheter " när han talade till sina 142 miljoner följare , bara timmar efter det att kraven rapporterades .
" Nej nej nej nej nej .
Vad de sa idag var falska nyheter " , sa den femfaldiga Ballon d ' Or @-@ vinnaren till kameran .
" De vill marknadsföra sig genom att använda mitt namn .
Det är normalt .
De vill bli kända genom att använda mitt namn , men det är en del av jobbet .
Jag är en lycklig man och allt bra " , sa spelaren och log .
Ronaldos advokater förbereder sig för att stämma Der Spiegel över påståenden , som de har kallat " en otillåtet rapportering av misstankar om integritet " , enligt Reuters .
Advokat Christian Schertz sa att spelaren skulle söka ersättning för " moralskada till ett belopp som motsvarar överträdelsens allvar , vilket förmodligen är en av de mest allvarliga kränkningarna av personliga rättigheter de senaste åren " .
Den påstådda händelsen sägs ha ägt rum i juni 2009 i en svit på Palms Hotel and Casino i Las Vegas .
Efter att ha träffats på en nattklubb gick Ronaldo och Mayorga tillbaka till spelarens rum , där han enligt uppgift ska ha våldtagit henne analt , enligt handlingar inlämnade vid Clark County District Court i Nevada .
Mayorga hävdar att Ronaldo föll på knä efter den påstådda händelsen och berättade för henne att han var " 99 procent " en " bra kille " sviken av den " sista procenten " .
Enligt dokumenten hade Ronaldo bekräftat att paret hade sex , men att det var med samtycke .
Mayorga hävdar också att hon gick till polisen och tog fotografier av sina skador på ett sjukhus , men kom senare överens om en förlikning eftersom hon kände sig " rädd för vedergällning " och var orolig för att " bli förödmjukad offentligt " .
34 @-@ åringen säger att hon nu försöker upphäva förlikningen eftersom hon fortsätter att traumatiseras av den påstådda händelsen .
Ronaldo var på väg att gå med i Real Madrid från Manchester United vid tiden för det påstådda överfallet , och i sommar flyttade han till den italienska jätten Juve i en överenskommelse på100 miljoner euro .
Brexit : Storbritannien " kommer för alltid ångra " att förlora biltillverkare
Storbritannien " skulle ångra det för alltid " om man förlorade sin status som världsledande inom biltillverkning efter Brexit , har affärsminister Greg Clark sagt .
Han tillade att det var " oroande " att Toyota UK hade berättat för BBC att om Storbritannien lämnade EU utan en överenskommelse kommer de att tillfälligt upphöra med produktionen vid fabriken i Burnaston , nära Derby .
" Vi behöver en överenskommelse " sade Clark .
Den japanska bilproducenten meddelade att effekterna av förseningar vid gränsen i händelse av att inget avtal sluts skulle kunna resultera i förlorade jobb .
Burnaston @-@ fabriken - som tillverkar Toyota ' s Auris och Avensis - producerade nästan 150 000 bilar i fjol , varav 90 % exporterades till resten av EU .
" Min åsikt är att om Storbritannien lämnar EU i slutet av mars kommer vi att se produktionsstopp i vår fabrik " , säger Marvin Cooke , Toyotas vd på Burnaston .
Andra brittiska biltillverkare har kommunicerat sin oro om att lämna EU utan en överenskommelse om hur gränsöverskridande handel kommer att fungera , inklusive Honda , BMW och Jaguar Land Rover .
BMW säger till exempel att det kommer att stänga sin Mini @-@ anläggning i Oxford i en månad efter Brexit .
Huvudproblemen gäller vad bilproducenterna säger är risker för försörjningskedjan i händelse av en Brexit utan uppgörelse .
Toyotas produktionslinje drivs på " just @-@ in @-@ time " -basis , med delar som kommer var 37:e minut från leverantörer i både Storbritannien och EU för bilar som beställts .
Om Storbritannien lämnar EU utan en överenskommelse den 29 mars kan det leda till störningar vid gränsen som branschen säger kan leda till förseningar och brist på delar .
Det skulle vara omöjligt för Toyota att hålla mer än en dags förbrukning i lager på dess Derbyshire @-@ fabrik , sa företaget , och därav skulle produktionen tvingas stoppas .
Clark sa att Theresa May ' s Chequers plan för framtida förbindelser med EU är " exakt kalibrerad för att undvika kontroller vid gränsen " .
" Vi behöver en uppgörelse . Vi vill ha den bästa överenskommelsen som möjliggör , som jag säger , inte bara framgång för närvarande att uppskattas nu , men för oss att ta tag i denna möjlighet " . sa han till BBC Radio 4:s program Today .
" Utsagorna från inte bara Toyota men andra tillverkare är att vi absolut måste kunna fortsätta det som har varit en mycket framgångsrik uppsättning av leverantörskedjor " .
Toyota kunde inte säga hur länge produktionen skulle stoppas , men på längre sikt varnade för att ökade kostnader skulle minska anläggningens konkurrenskraft och så småningom kosta jobb .
Peter Tsouvallaris , som har arbetat i Burnaston i 24 år och är ledare för Unite @-@ fackföreningen vid fabriken , sa att hans medlemmar är alltmer oroliga : " Min erfarenhet är att dessa jobb aldrig kommer tillbaka .
En regeringstjänsteman sa : " Vi har lagt fram en exakt och trovärdig plan för vårt framtida förhållande till EU " .
Trumps möte med Rosenstein kan försenas igen , säger Vita huset
Donald Trumps möte med biträdande justitieminister Rod Rosenstein skulle kunna " skjutas på ännu en vecka " medan kampen mot den till högsta domstolen nominerade Brett Kavanaugh fortsätter , sade Vita huset på söndagen .
Rosenstein övervakar arbetet med specialrådgivaren Robert Mueller , som undersöker rysk inblandning i valet , förbindelser mellan Trump och Ryssland och presidentens potentiella hindrande för rättvisa .
Huruvida Trump kommer att sparka den biträdande justitieministern , och därigenom äventyra Muellers självständighet , har gett bränsle åt Washingtonskvaller i månader .
Tidigare denna månad rapporterade New York Times att Rosenstein diskuterade möjligheten att bära avlyssningsutrustning för att spela in konversationer med Trump samt möjligheten att avsätta presidenten via det 25:e tillägget av den amerikanska konstitutionen .
Rosenstein förnekade rapporten .
Men i måndags gick han till Vita huset , och rapporter om att han skulle avgå framkom .
Istället tillkännagavs ett möte med Trump , som då var i FN:s högkvarter i New York , som ska hållas på torsdagen .
Trump sa att han skulle " föredra " att inte sparka Rosenstein men sedan blev mötet försenat för att undvika en konflikt med senatens juridiska utskotts förhör där Kavanaugh och en av de kvinnor som har anklagat honom för sexuell oegentlighet , Dr Christine Blasey Ford , båda vittnade .
På fredagen ​ ​ beställde Trump en en @-@ veckas FBI @-@ undersökning av anklagelser mot Kavanaugh , vilket ytterligare försenade en full omröstning i senaten .
Trumps pressekreterare , Sarah Sanders , talade i Fox News på söndagen .
När hon tillfrågades om mötet med Rosenstein sa hon : " Ett datum för det har inte fastställts , det kan ske den här veckan , eller en senareläggning med en vecka med tanke på alla andra saker som händer vid högsta domstolen .
Men vi får se , och jag gillar alltid att hålla pressen uppdaterad . "
Vissa reportrar skulle bestrida det påståendet : Sanders har inte haft en presskonferens från Vita huset sedan den 10 september .
Värden Chris Wallace frågade varför .
Sanders sa att bristen på presskonferenser inte berodde på något ogillande gentemot TV @-@ reportrar som " spelar för galleriet " , även om hon sa : " Jag håller med om det faktum att de spelar för galleriet " .
Hon sa sedan att direktkontakt mellan Trump och pressen kommer att öka .
" Presidenten håller flera frågesessioner än någon president före honom " , sa hon och tillade utan att citera bevis : " Vi har tittat på dessa siffror " .
Konferenser kommer fortfarande att äga rum , sade Sanders , men " om pressen får chansen att ställa frågor direkt till USA:s president är det oändligt mycket bättre än att prata med mig .
Vi försöker att göra detta ofta och ni har sett oss göra mycket under de senaste veckorna och det kommer ersätta presskonferenser , och ni kan då ställa frågor direkt till USA : s president " .
Trump svarar regelbundet på frågor när han lämnar Vita huset eller deltar i öppna sessioner eller presskonferenser med besökande dignitärer .
Solo @-@ presskonferenser är sällsynta .
I New York den här veckan visade presidenten kanske varför , med spontana uttalanden och ibland bisarra framträdanden inför de samlade reportrarna .
Hälsosminister skriver till medarbetare från EU vid NHS Skottland med hänsyn till oro om Brexit
Hälsoministern har skrivit till EU @-@ personal som arbetar i Skottlands NHS för att uttrycka landets tacksamhet och önskan att de ska stanna kvar efter Brexit .
Jeane Freeman , MSP , skickade ett brev mindre än sex månader innan Storbritannien drar sig ur EU .
Den skotska regeringen har redan åtagit sig att täcka kostnaden för avvecklade statusansökningar för EU @-@ medborgare som arbetar i landets decentraliserade offentliga sektor .
I brevet skrev Freeman : " Under sommaren har förhandlingarna mellan Storbritannien och EU om utträde fortsatt , inför beslut som förväntas komma i höst .
Men den brittiska regeringen har också intensifierat sina förberedelser inför ett eventuellt scenario utan överenskommelse .
Jag vet att detta måste vara en mycket oroande tid för er alla .
Därför vill jag upprepa hur mycket jag värderar varje medarbetares insats , oavsett nationalitet .
Kollegor från hela EU , och resten av världen , ger värdefull erfarenhet och kompetens som stärker och förbättrar hälsovårdens arbete och gynnar de patienter och samhällen vi tjänar .
Skottland är definitivt ditt hem och vi vill verkligen att du ska stanna här " .
Christion Abercrombie genomgår akut kirurgi efter att han drabbats av huvudskada
Tennessee State Tigers linjeback Christion Abercrombie genomgick en akut operation efter att ha drabbats av en huvudskada i lördagens förlust med 31 @-@ 27 mot Vanderbilt Commodores , rapporterade Tennesseans Mike Organ .
Tennessee States huvudtränare Rod Reed berättade för reportrarna att skadan skedde strax före halvtid .
" Han kom till sidlinjen och bara kollapsade " , sade Reed .
Tränare och medicinsk personal gav Abercrombie syre på sidolinjen innan han placerades på en bår fördes ut för vidare utvärdering .
En representant från Tennessee State berättade för Chris Harris från WSMV i Nashville , Tennessee , att Abercrombie opererades vid sjukhuset Vanderbilt Medical Center .
Harris tillade att " det finns inga uppgifter om typen / omfattningen av skadan än " och Tennessee State försöker ta reda på när skadan inträffade .
Abercrombie , en redshirt andraårsstudent , är i sin första säsong med Tennessee State efter en överföring från Illinois .
Han hade totalt fem tacklar på lördagen innan han lämnade matchen , vilket gav honom en säsongtotal på 18 tacklar .
Utländska köpare kommer att debiteras högre stämpelskatt när de köper en fastighet i Storbritannien
Utländska köpare får betala högre stämpelskatt när de köper egendom i Storbritannien , och de extra pengarna används för att hjälpa hemlösa , enligt Tory @-@ partiets nya planer
Åtgärden ska neutralisera Corbyns framgångar med att attrahera unga väljare
Höjningen av stämpelskatten kommer att gälla dem som inte betalar skatt i Storbritannien
Det brittiska finansdepartementet räknar med att få in upp till 120 miljoner pund om året för att hjälpa de hemlösa
Utländska köpare ska få betala en högre stämpelskatt när de köper egendom i Storbritannien . De extra pengarna ska användas för att hjälpa hemlösa , vilket kommer att tillkännages av premiärminister Theresa May i dag .
Åtgärden kommer att uppfattas som ett försök att neutralisera Jeremy Corbyns framgångar med att attrahera unga väljare med löften om bostäder med mer överkomliga priser och att sikta in sig på höginkomsttagare .
Höjningen av stämpelskatten kommer att tas ut av individer och bolag som inte betalar skatt i Storbritannien . Extrapengarna ska ge en skjuts åt regeringens satsning på att bekämpa hemlösheten .
Den extra avgiften tillkommer utöver den nuvarande stämpelskatten , inklusive de högre nivåerna som infördes för två år sedan på fritidsbostäder och bostäder som köps för att hyras ut . Den kan komma att ligga på upp till tre procent .
Finansdepartementet tror att åtgärden kommer att dra in upp till 120 miljoner pund per år .
Uppskattningsvis 13 procent av de nybyggda fastigheterna i London köps av personer som bor utanför Storbritannien . Detta driver upp priserna och gör det svårare för förstagångsköpare att få in en fot på bostadsmarknaden .
Många välbärgade områden i landet , särskilt i huvudstaden , har blivit spökstäder på grund av det höga antalet utländska köpare som tillbringar större delen av sin tid utomlands .
Det nya utspelet kommer bara några veckor efter det att Boris Johnson efterfrågade en minskning av stämpelskatten för att hjälpa fler unga att kunna köpa sin första bostad .
Han anklagade stora byggbolag för att hålla priserna uppe genom att köpa upp mark utan att använda den , och uppmanade Theresa May att avstå från kvoter på bostäder med överkomliga priser för att lösa Storbritanniens " bedrövliga bostadssituation " .
Jeremy Corbyn har lanserat en uppseendeväckande räcka förslag till bostadsreformer , däribland hyrestak och ett slut på vräkningar utan hyresgästens förskyllan .
Han vill också ge kommunerna större möjlighet att bygga nya bostäder .
Theresa May säger : " Förra året sade jag att jag skulle ägna min tid som premiärminister åt att återupprätta den brittiska drömmen , att livet ska bli bättre för varje ny generation .
Det innebär att lösa problemen på bostadsmarknaden .
Storbritannien kommer alltid att vara öppet för människor som vill bo , arbeta och bygga upp ett liv här .
Men det kan inte stå rätt till när det är lika lätt för personer som inte bor i Storbritannien , och även för företag som är baserade i utlandet , att köpa bostäder som för hårt arbetande invånare i vårt land .
Drömmen om att äga sin bostad har för alltför många människor blivit just en avlägsen dröm , och hemlösheten är fortfarande ett ovärdigt faktum " .
Jack Ross : " Mitt slutliga mål är att träna Skottland "
Sunderland @-@ ledaren Jack Ross säger att hans " slutliga mål " är att någon gång bli Skottlands tränare .
Den 42 @-@ årige skotten ser fram emot utmaningen att blåsa liv i klubben från nordöstra England , som för närvarande ligger på tredje plats i League One , tre poäng från toppen .
Han flyttade till Stadium of Light i somras efter att ha lett St Mirren tillbaka till Scottish Premiership förra säsongen .
" Jag ville spela för mitt land som spelare .
Jag spelade en match i B @-@ landslaget och det var allt " , säger Ross till BBC Scotlands Sportsound .
" Men när jag växte upp tittade jag mycket på Skottland på Hampden med min pappa , och det har alltid lockat mig tillbaka .
Men den chansen kan bara komma om jag lyckas med att leda en klubb " .
Bland Ross företrädare som tränare för Sunderland finns Dick Advocaat , David Moyes , Sam Allardyce , Martin O ' Neill , Roy Keane , Gus Poyet och Paulo Di Canio .
Den tidigare ledaren för Alloa Athletic säger att han inte var orolig för att efterträda så etablerade namn i en så stor klubb . Han har tidigare tackat nej till erbjudanden från Barnsley och Ipswich Town .
" Just nu bedömer jag framgång utifrån svaret på frågan " kan jag få den här klubben tillbaka till Premier League ? "
Den här klubben hör absolut hemma i Premier League , med tanke på dess struktur och talanger " , säger han .
" Det är inte lätt att komma dit , men jag skulle nog bara se mig själv som framgångsrik här om jag kan få klubben tillbaka dit " .
Ross har bara varit tränare i tre år , efter en period som assisterande tränare i Dumbarton och en 15 månader lång sejour som medlem av Hearts tränarteam .
Då hjälpte han Alloa att komma tillbaka från nedflyttning till tredje divisionen , och lyfte St Mirren från att vara nära nedflyttning till att bli vinnare av mästerskapstiteln säsongen därpå .
Ross säger att han är mer tillfreds nu än någonsin under sin spelarkarriär i Clyde , Hartlepool , Falkirk , St Mirren och Hamilton Academical .
" Det var antagligen ett vägskäl " , minns han och syftar på när han tog befälet över Alloa .
" Jag trodde verkligen att ledarskap var helt rätt för mig , på ett helt annat sätt än att spela .
Det låter konstigt , för jag hade okej resultat och kunde leva hyfsat på det . Dessutom hade jag vissa stora framgångar .
Men att spela kan vara tufft .
Det är mycket man måste ta sig igenom varje vecka .
Det är fortfarande stress och press på jobbet för mig , men att träna känns helt rätt .
Jag har alltid velat träna och nu gör jag det . Jag mår bättre än jag har gjort någonsin under hela mitt vuxna liv " .
Lyssna på hela intervjun i Sportsound , söndagen den 30 september på Radio Scotland mellan 12 : 00 och 13 : 00
En undersökning visar att den perfekta tiden att ta en öl är 17 : 30 på en lördag
Sommarens värmebölja har inneburit ökade intäkter för landets kämpande pubar , men restaurangkedjorna har fått större press på sig .
Siffror visade att pub- och barkoncerner ökade försäljningen med 2,7 % i juli , men restaurangernas intäkter sjönk med 4,8 % .
Peter Martin från företagsrådgivningsbolaget CGA , som har sammanställt siffrorna , sade : " Fortsatt vackert väder och det faktum att England blev kvar i VM längre än väntat innebar att vi fick se ett liknande mönster i juli jämfört med juni , då pubarna gick upp med 2,8 % . Restaurangerna fick dock ännu större svårigheter .
Minskningen i restaurangernas omsättning med 1,8 % i juni blev bara värre i juli .
Pubar och barer som framför allt erbjuder drycker uppvisade det absolut bästa resultatet med siffror för samma period förra året som hade gått upp mer än restaurangerna hade gått ner .
Pubar som erbjuder mat hade det också svårt i det vackra vädret , även om det inte var lika dramatiskt som för restaurangägare .
Folk verkar bara ha velat gå ut och dricka något .
Utslaget på förvaltade pubar och barer gick dryckesförsäljningen upp med 6,6 % den månaden , och matförsäljningen ner med 3 % " .
Paul Newman på serverings- och nöjesbranschanalytikern RSM säger : " De här resultaten är en fortsättning på tendensen vi har sett sedan slutet av april .
Vädret och stora sportevenemang är fortfarande de viktigaste faktorerna när det gäller försäljning på storköksmarknaden .
Det är ingen överraskning att restaurangkoncernerna fortfarande har svårigheter , även om en försäljningsminskning på 4,8 % varje år är särskilt svårt att hantera utöver pågående kostnadstryck .
Den långa varma sommaren kunde inte ha kommit mer olägligt för företag som drivs av matförsäljning . Tiden får utvisa om de mer måttliga temperaturerna som vi har haft i augusti ger någon välbehövd respit " .
Den totala försäljningsökningen utslaget på pubar och restauranger , inklusive nyöppnade inrättningar , låg på 2,7 % i juli . Det återspeglar det faktum att det nu lanseras färre nya varumärken .
Branschförsäljningsövervakaren Coffer Peach Tracker för pub- bar- och restaurangbranschen i Storbritannien samlar in och analyserar uppgifter om hur det går för 47 aktiva koncerner med en sammanlagd omsättning på över 9 miljarder pund , och är ett etablerat riktmärke i branschen .
Ett av fem barn har hemliga konton på sociala medier som de döljer för sina föräldrar
En undersökning visar att ett av fem barn , ibland så unga som 11 år , har hemliga konton på sociala medier som de döljer för sina föräldrar och lärare
En undersökning bland 20 000 elever på högstadiet och gymnasiet visar en ökning av antalet falska Instagramsidor
Resultatet har ökat oron för att det är sexuellt innehåll som läggs upp där
20 % av eleverna uppgav att de hade ett " huvudkonto " som de visade för sina föräldrar
Ett av fem barn , vissa så unga som 11 år , skapar konton på sociala medier som de håller hemliga för vuxna .
En undersökning bland 20 000 elever i högstadiet och gymnasiet visade en snabb ökning av antalet " falska Instakonton " , en hänvisning till bilddelningstjänsten Instagram .
Resultatet har spätt på oron för att det är sexuellt innehåll som postas där .
20 % av eleverna uppgav att de har ett städat " huvudkonto " som de kan visa för sina föräldrar , och så har de även privata konton .
En mamma som snubblade över hennes 13 @-@ åriga dotters hemliga sida hittade en tonåring som uppmanade andra att " våldta mig " .
Enligt studien , som utfördes av organisationerna Digital Awareness UK och Headmasters och Headmistresses Conference ( HMC ) of independent schools , hade 40 % av barnen mellan 11 och 18 år två profiler , och hälften av dem erkände att de hade privata konton .
Ordföranden för HMC , Mike Buchanan , säger : " Det är oroande att så många tonåringar lockas att skapa platser på internet där föräldrar och lärare inte hittar dem " .
Eilidh Doyle kommer att vara " idrottarnas röst " i styrelsen för det skotska friidrottsförbundet , Scottish Athletics
Eilidh Doyle har blivit invald i styrelsen för Scottish Athletics som extern styrelsemedlem vid det styrande organets årsstämma .
Doyle är Skottlands mest prisade friidrottare , och ordföranden Ian Beattie beskriver valet som en enastående möjlighet för dem som leder idrotten att dra nytta av hennes breda erfarenhet på internationell nivå det senaste decenniet .
" Eilidh har vunnit stor respekt i hela den skotska , brittiska och internationella idrottsvärlden , och vi är säkra på att idrottarna i Skottland skulle ha stor nytta av att hon blir en medlem av styrelsen " , säger Beattie .
Doyle säger : " Jag vill gärna vara en röst för idrottarna och jag hoppas att jag kan bidra och hjälpa till att leda sporten i Skottland " .
Amerikanen , som vann 200 meter och 400 meter vid OS i Atlanta 1996 , har totalt fyra olympiska guld och är nu expertkommentator på BBC . Han förlorade förmågan att gå efter en mini @-@ stroke .
Han skriver på Twitter : " I dag för en månad sedan fick jag en stroke .
Jag kunde inte gå .
Läkarna sade att tiden fick utvisa om jag skulle återhämta mig , och i vilken utsträckning .
Det har varit hårt arbete , men jag har återhämtat mig helt och hållet , lärt mig gå igen och nu gör jag rörlighetsövningar !
Tack för all uppmuntran ! "
Reklam för bröstpumpar som jämför mammor med kor delar internet
Ett företag som säljer bröstpumpar har orsakat meningsskiljaktigheter på internet med en annons som jämför ammande mammor med kor som blir mjölkade .
För att uppmärksamma lanseringen av vad som sägs vara " världens första tysta bärbara bröstpump " har konsumentteknikbolaget Elvie släppt en musikvideoinspirerad reklamfilm med humoristiskt anslag för att visa på vilken frihet den nya pumpen ger mammor som pumpar bröstmjölk .
Fyra verkliga mammor dansar i en höfylld lada med kor till en låt med textrader som : " Ja , jag mjölkar mig själv , men har ingen svans " och " Om du inte visste det , så är det här inget juver , utan tuttar " .
Refrängen fortsätter : " Pumpa ut , pumpa ut , jag matar bebisarna , pumpa ut , pumpa ut , jag mjölkar damerna " .
Men reklamfilmen , som har publicerats på företagets Facebook @-@ sida , har orsakat strid på internet .
Filmen har fått 77 000 visningar och hundratals kommentarer , och har mött blandade reaktioner från tittarna . Många säger att den kastar ljus över mejeriindustrins " fasor " .
" Ett mycket dåligt beslut att använda kor för att marknadsföra den här produkten .
Precis som vi måste de bli gravida och föda för att kunna producera mjölk , men deras ungar tas ifrån dem bara några dagar efter födseln " , skriver en person .
Elvie bröstpump kan bäras diskret i en amningsbehå ( Elvie / Mother )
En annan kommenterar : " Man förstår att det är traumatiskt för både mamma och barn .
Men visst , varför inte använda dem för att göra reklam för en bröstpump för mödrar som får behålla sina barn ? "
Ytterligare någon tillägger : " Vilken verklighetsfrånvänd reklamfilm . "
Andra försvarar filmen , och en kvinna medger att hon tycker att sången är " hysteriskt rolig " .
" Jag tycker att det här är genialiskt .
Jag skulle ha skaffat en om jag fortfarande ammade .
Att pumpa fick mig att känna mig precis som en ko .
Reklamfilmen är lite galen , men jag tog den för vad den var .
Det här är en genialisk produkt " , skriver någon .
En annan kommenterar : " Det här är en rolig reklamfilm som vänder sig till mammor som pumpar ( ofta på arbetsplatsen eller på toaletten ) och känner sig som " kossor " " .
Det här är inte en film som hyllar eller fördömer mejeriindustrin " .
I slutet av filmen avslöjar kvinnorna att de alla har dansat med den diskreta pumpen instoppad i behån .
Konceptet bakom kampanjen är baserat på att många kvinnor som pumpar mjölk säger att de känner sig som kor .
Men Elvie @-@ pumpen är helt tyst , har inga kablar eller rör och kan bäras diskret i en amningsbehå , vilket ger kvinnorna frihet att röra sig , hålla sina bebisar och till och med gå ut medan de pumpar .
Ana Balarin är delägare och ECD på Mother , och hon säger : " Elvie @-@ pumpen är en så revolutionerande produkt att den förtjänar en djärv och provokativ lansering .
Genom att dra en parallell mellan kvinnor som pumpar bröstmjölk och mjölkkor ville vi sätta ljus på bröstpumpning och utmaningarna med det , samtidigt som vi på ett underhållande och lätt igenkännbart sätt visar vilken otrolig frihetskänsla den nya pumpen ger .
Det här är inte första gången Elvie @-@ pumpen skapar rubriker .
Under Londons modevecka framträdde en tvåbarnsmamma på catwalken med kläder av designern Marta Jakubowski samtidigt som hon använde produkten .
Hundratals migrantbarn flyttade i tysthet till ett tältläger nära gränsen i Texas
Antalet frihetsberövade migrantbarn har skjutit i höjden även om antalet personer som korsar gränsen varje månad är relativt oförändrat . Detta beror delvis på att hätsk retorik och hård politik som har införts av regeringen Trump har gjort det svårare att placera barnen hos referenspersoner .
Tidigare har de flesta referenspersoner själva varit papperslösa invandrare , och rädda att sätta sina egna möjligheter att stanna i landet på spel genom att förklara sig villiga att ta emot ett barn .
Risken ökade i juni när federala myndigheter tillkännagav att potentiella referenspersoner och andra vuxna medlemmar i hushållet skulle vara tvungna att lämna fingeravtryck , och att uppgifterna skulle delas med invandringsmyndigheterna .
Förra veckan vittnade Matthew Albence , en högre tjänsteman på Invandrings- och tullmyndigheten , inför kongressen om att myndigheten hade gripit dussintals personer som hade ansökt om att få vara referenspersoner åt ensamkommande minderåriga .
Myndigheten bekräftade senare att 70 % av dem som greps inte var kända av brottsbekämpande myndigheter sedan tidigare .
" Nästan 80 % av de personer som antingen själva är referenspersoner eller familjemedlemmar till referenspersoner befinner sig olagligt i landet , och en stor del av dem är kriminella utlänningar .
Så vi fortsätter att förfölja dessa individer " , sade Albence .
För att hantera barnens ärenden snabbare har tjänstemän infört nya regler som kräver att vissa av dem ska infinna sig i rätten inom en månad efter de att de frihetsberövades , snarare än efter 60 dagar , vilket tidigare var praxis , enligt personal på förläggningarna .
Många av dem är närvarande på videolänk snarare än personligen för att föra sin talan för rättslig status inför en invandringsdomare .
De som inte bedöms ha rätt till skydd deporteras snabbt .
Ju längre barn är frihetsberövade desto mer sannolikt är det att de drabbas av ångest eller depression , vilket kan leda till våldsamma utbrott eller flyktförsök , enligt personal på förläggningarna och rapporter som har kommit från systemet de senaste månaderna .
Förespråkare säger att oron stiger vid större anläggningar som Tornillo , där tecken på att ett barn har det svårt mer sannolikt ignoreras , på grund av anläggningens storlek .
De tillägger att om barn flyttas till tältstaden utan att få tillräckligt med tid att förbereda sig känslomässigt och ta farväl av vänner kan förvärra de trauman många redan brottas med .
Syrien kräver att amerikanska , franska och turkiska " ockupationsstyrkor " ska dra sig tillbaka omedelbart
I ett tal till FN:s generalförsamling uppmanade utrikesminister Walid al @-@ Moualem också syriska flyktingar att komma hem igen , trots att kriget i landet är inne på sitt åttonde år .
Moualem , som också är vice premiärminister , sade att de utländska styrkorna befinner sig illegalt på syrisk mark , under förevändningen att bekämpa terrorism , och " kommer att hanteras i enlighet med detta " .
" De måste dra sig tillbaka omedelbart och villkorslöst " , sade han till generalförsamlingen .
Moualem underströk att " kriget mot terrorn är nästan över " i Syrien , där fler än 360 000 människor har dött sedan 2011 , och miljoner lämnat sina hem .
Han sade att regeringen i Damaskus skulle fortsätta att " utkämpa detta heliga slag tills vi har befriat alla syriska territorier " både från terrorgrupper och " all olaglig utländsk närvaro " .
USA har ungefär 2 000 soldater i Syrien , som främst utbildar och ger råd åt både kurdiska styrkor och syriska araber som är motståndare till president Bashar al @-@ Assad .
Frankrike har mer än 1 000 soldater på marken i det krigshärjade landet .
Vad gäller flyktingarna sade Moualem att det omständigheterna är goda för att de ska komma hem , och anklagade " vissa västländer " för att " sprida irrationell rädsla " som förmår flyktingar att hålla sig borta .
" Vi har uppmanat det internationella samfundet och humanitära organisationer att underlätta deras återvändande " , sade han .
" De politiserar något som borde vara en rent humanitär fråga " .
USA och EU har varnat för att det inte blir någon hjälp till återuppbyggnad till Syrien förrän det finns en politisk överenskommelse mellan Assad och oppositionen att avsluta kriget .
FN @-@ diplomater säger att en färsk överenskommelse mellan Ryssland och Turkiet att upprätta en buffertzon i det sista stora rebellfästet Idlib har skapat en möjlighet att gå vidare med politiska samtal .
Det rysk @-@ turkiska avtalet avstyrde ett storskaligt anfall av ryskstödda syriska trupper mot provinsen , som har tre miljoner invånare .
Moualem betonade dock att överenskommelsen hade " tydliga deadlines " , och uttryckte hopp om att ett militärt ingripande skulle riktas mot jihadister , inklusive krigare från den Al Qaida @-@ kopplade Nusrafronten , som " kommer att utplånas " .
FN @-@ sändebudet Staffan de Mistura hoppas snart kunna sammankalla de första mötena i en ny kommitté som består av regeringsmedlemmar och medlemmar av oppositionen , för att göra ett utkast till efterkrigskonstitution för Syrien och bana väg för val .
Moualem ställde upp villkor för den syriska regeringens deltagande i kommittén och sade att gruppens arbete skulle begränsas till " översyn av artiklarna i den nuvarande konstitutionen " , och varnade för inblandning .
Varför Donald Trump kommer att vinna ett omval
Med den logiken skulle Donald Trump vinna omvalet 2020 om inte hans presidentskap avslutas i förtid genom riksrätt och skandal , vilket många liberala tittare troligen hoppas på .
I det som utan tvivel skulle vara " den mest dramatiska finalen på ett presidentskap någonsin ! "
I nuläget finns inga tecken på att tittarna har tröttnat .
Sedan 2014 har tittarsiffrorna på bästa sändningstid mer än fördubblats till 1,05 miljoner på CNN , och är nästan tre gånger så höga , 1,6 miljoner , på MSNBC .
Fox News har ett genomsnitt på 2,4 miljoner tittare på bästa sändningstid , vilket är en ökning från 1,7 miljoner för fyra år sedan , enligt Nielsen . MSNBC:s " The Rachel Maddow Show " har toppat listorna för kabelkanaler med så många som 3,5 miljoner tittare under stora nyhetskvällar .
" Det här är som en eld som folk dras till , för det är något vi inte förstår " , sade Neal Baer , som driver showen för ABC:s drama " Designated Survivor " , som handlar om en kabinettssekreterare som blir president efter att en attack har förstört Capitolium .
Nell Scovell är mångårig komediförfattare och har skrivit " Just the Funny Parts : And a Few Hard Truths About Sneaking Into the Hollywood Boys " Club " . Hon har en annan teori .
Hon minns en taxifärd i Boston före valet 2016 .
Föraren berättade att han skulle rösta på Donald Trump .
Varför då ? frågade hon .
" Han sade , " För att han får mig att skratta " " , berättar Nell Scovell för mig .
I kaoset finns ett underhållningsvärde .
Givetvis är det så att till skillnad från allt annat på TV , så kan rapporteringen från Washington avgöra framtiden för rättsfallet i abortfrågan , Roe vs Wade , huruvida invandrarfamiljer kan återförenas och den globala ekonomins välmående .
Att stänga av är en lyx som bara de mest privilegierade tittarna har råd med .
Ändå går det utöver att vara en informerad medborgare när man plötsligt har suttit och tittat i sex timmar på en expertpanel som debatterar Bob Woodwards användande av " djupa bakgrundskällor " till sin bok " Fear " , Paul Manaforts bomberjacka av strutsläder för 15 000 dollar ( " ett plagg fyllt av hybris " , som Washington Post sa ) och innebörden i Stormy Daniels makabra beskrivningar av Donald Trumps , hm , anatomi .
Jag kommer själv aldrig att se på Super Mario på samma sätt igen .
" En del av det han gör som får det att kännas som en realityserie är att han kommer med något varje kväll " , sade Brent Montgomery , vd för Wheelhouse Entertainment och skapare av " Pawn Stars " , om Trump @-@ följetongens roterande rollbesättning och dagliga intriger ( mucka gräl med NFL , lovorda Kim Jong @-@ un ) .
Om man missar ett enda avsnitt hamnar man på efterkälken .
När jag talade med tv @-@ producenten mr Fleiss den här veckan var det sol och 27 grader utanför hans hus på norra Kauai på Hawaii , men han satt och ugglade inomhus och tittade på MSNBC samtidigt som han spelade in en sändning från CNN .
Han kunde inte slita sig , inte när Brett Kavanaugh skulle ställas inför senatens justitieutskott och Högsta Domstolens framtid låg i vågskålen .
" Jag kommer ihåg när vi gjorde alla de där galna programmen förr i tiden och folk sade : " Det här är början till slutet på den västliga civilisationen " " , sade mr Fleiss till mig .
" Jag trodde att det var någon sorts skämt , men det visade sig att de hade rätt " .
Amy Chozick , som är fristående skribent för The Times och skriver om ekonomi , politik och media , är författare till biografin " Chasing Hillary " .
Pengar utifrån strömmar in i den jämnaste kapplöpningen någonsin inför mellanårsvalet
Det är inte förvånande att Pennsylvanias 17:e kongressdistrikt tar emot massor av pengar . Det är tack vare en omstrukturering av ett kongressdistrikt som har gjort att två ledamöter nu tävlar om samma plats .
Detta nyligen omritade förortsdistrikt i Pittsburg representeras av demokraten Conor Lamb , som fick sin plats i ett annat distrikt vid ett specialval förra våren .
Lamb kampanjar mot en annan ledamot , republikanen Keith Rothfus . Han representerar för närvarande det gamla 12:e distriktet i Pennsylvania , som i stor utsträckning överlappar det nya 17:e distriktet .
Kartorna ritades om efter det att Pennsylvanias Högsta Domstol i januari beslutade att de gamla distrikten var konstitutionsvidrigt ändrade till republikanernas fördel .
Kapplöpningen i det nya 17:e distriktet har orsakat en kampanjfinansieringsstrid mellan de största partiernas ekonomisektioner , Democratic Campaign Congressional Committee , ( DCCC ) och National Republican Campaign Committee ( NRCC ) .
Lamb blev ett bekant namn i Pennsylvania efter en knapp vinst i ett brett bevakat specialval i mars till Pennsylvanias 18:e kongressdistrikt .
Den platsen hade innehafts av en republikan i över ett decennium , och president Donald Trump vann distriktet med 20 poäng .
Politiska experter hade gett demokraterna ett visst försprång .
USA övervägde att bestraffa El Salvador för Kinastöd men backade sedan
Diplomater noterade att Dominikanska republiken och Panama redan hade erkänt Peking , med lite motstånd från Washington .
Donald Trump hade ett varmt möte med Panamas president Juan Carlos Varela i juni 2017 , och hade ett hotell i Panama , tills delägarna vräkte Trumporganisationens ledarteam .
Tjänstemän på det amerikanska utrikesdepartementet beslutade att kalla hem cheferna för de amerikanska beskickningarna i El Salvador , Dominikanska republiken och Panama på grund av " nyss fattade beslut att inte längre erkänna Taiwan " , sade departementets talesperson Heather Nauert i ett uttalande tidigare den här månaden .
Men man planerade bara sanktioner mot El Salvador , som fick uppskattningsvis 140 miljoner dollar i amerikanskt bistånd 2017 . Pengarna skulle bland annat gå till narkotikakontroll och utveckling och utgöra ekonomiskt stöd .
De föreslagna sanktionerna , däribland minskat ekonomiskt bistånd och riktade visumrestriktioner , skulle ha slagit hårt mot det centralamerikanska landet med dess höga arbetslöshet och mordstatistik .
Samtidigt som de interna mötena fortskred sköt amerikanska och centralamerikanska tjänstemän upp en högnivåkonferens med fokus på säkerhet och ekonomiskt välstånd för att följa upp ett liknande möte förra året , som sågs som ett steg i rätt riktning för att hindra migranter från att bege sig till USA .
Men i mitten av september gjorde höga tjänstemän inom administrationen klart att de ville att konferensen skulle äga rum , vilket i praktiken satte stopp för överväganden om sanktioner mot El Salvador .
Vicepresident Mike Pence ska nu tala på konferensen , som nu ska äga rum i mitten av oktober . Det är ett tecken på hur viktigt presidentadministrationen anser mötet vara , sade diplomaterna .
Och de tre amerikanska sändebuden återvände i tysthet till El Salvador , Panama och Dominikanska republiken utan några nya hårda budskap eller bestraffningar från Washington .
En talesperson för John Bolton från Vita Huset avböjde att kommentera detaljerna i debatten , vilka beskrevs av de tre amerikanska tjänstemännen , varav två diplomater , som gick med på att diskutera de interna överläggningarna mot löfte om anonymitet .
Deras redogörelser bekräftades av en utomstående analytiker som står administrationen nära och som också uttalade sig anonymt .
Studera historien
Nästa oundvikliga steg kan bli den särskilde utredaren Robert Muellers rapport om Donald Trumps påstådda övergrepp i rättssak , som det nu finns påtagliga bevis för i offentliga register .
Mueller rapporteras också styra sin utredning mot huruvida Donald Trumps kampanj samarbetade med Ryssland i dess angrepp på det amerikanska valet .
Om kongressen skulle byta majoritet kommer Trump att hållas ansvarig inför den församlingen precis när han förbereder sig för att än en gång ställa upp i valet , och kanske slutligen inför en medborgarjury .
Det är många osäkra faktorer i detta , och jag vill inte påstå att Trump oundvikligen kommer att falla . Så inte heller hans kollegor i Europa .
Vi måste alla träffa olika val , på båda sidor av Atlanten , som kommer att påverka hur utdragen kampen kan bli .
1938 var tyska officerare redo att iscensätta en statskupp mot Hitler , om bara västländerna hade stått emot honom och ställt sig bakom tjeckoslovakerna i München .
Vi misslyckades , och missade ett tillfälle att undvika åren av blodbad som sedan följde .
Historien kretsar kring sådana avgörande händelser , och demokratins obevekliga frammarsch skyndas antingen på eller bromsas .
Amerikanerna står nu inför flera av dessa avgörande händelser .
Vad ska vi göra om Donald Trump ger biträdande justitieminister Rod Rosenstein , mannen som kontrollerar vad som ska hända med Muellers utredning , sparken ?
Rosenstein har varit i svårigheter ända sedan denna tidning rapporterade om att han förra året ska ha föreslagit att i hemlighet spela in presidenten , och spekulerat om att han inte skulle vara lämplig för ämbetet .
Rosenstein säger att The Times rapportering inte stämmer .
" Hur ska vi svara om den nyss begärda FBI @-@ utredningen av Brett Kavanaugh är ofullständig eller orättvis , eller om han får tillträda i Högsta Domstolen trots trovärdiga anklagelser om sexuella övergrepp och falskt vittnesmål ?
Och framför allt , kommer vi i mellanårsvalen att rösta på en kongress som håller Donald Trump ansvarig ?
Om vi misslyckas i dessa prövningar står demokratin inför en mörk period .
Men jag tror inte att vi kommer att misslyckas , på grund av den läxa jag lärde mig i Prag .
Min mamma var tjeckoslovakisk jude och deporterades till Auschwitz av samma nazistregim som en gång ockuperade mitt ambassadörsresidens .
Hon överlevde , invandrade till USA och 60 år senare skickade hon i väg mig för att tända sabbatsljus på det bord som var dekorerat med hakkorset .
Med det som arv , hur skulle jag kunna vara annat än optimist om framtiden ? "
Norman Eisen är mångårig medarbetare vid tankesmedjan Brookings Institution och ordförande i organisationen " Citizens for Responsibility and Ethics in Washington " , samt författare till " The Last Palace : Europe ' s Turbulent Century in Five Lives and One Legendary House " .
Graham Dorrans i Rangers är optimist inför mötet med Rapid Wien
Rangers tar emot Rapid Wien på torsdag . De vet att seger mot österrikarna efter den imponerande Spanienmatchen mot Villarreal som slutade oavgjort tidigare i månaden kommer att försätta dem i en stark ställning för att kvalificera sig från grupp G i Europa League .
En knäskada hindrade mittfältaren Graham Dorrans från att göra sitt första framträdande för säsongen , fram till 2 @-@ 2 @-@ matchen mot Villarreal . Men han tror att Rangers kan använda resultatet som en språngbräda mot större framgångar .
" Det var en bra poäng för oss , för Villarreal är ett bra lag " , säger 31 @-@ åringen .
" Vi gick in i matchen i tron att vi kunde få någonting , och gick därifrån med en poäng .
Vi kanske kunde ha fått in den i slutet , men i det stora hela var nog oavgjort ett rättvist resultat .
De var nog bättre i första halvlek . Vi kom igen i andra halvlek och var det bättre laget .
Nu på torsdag blir det en viktig kväll i Europa igen .
Förhoppningsvis kan vi få tre poäng , men det blir en tuff match . De fick ett bra resultat vid sin senaste match , men om vi har publiken med oss kan vi säkert rycka fram och få ett bra resultat .
Förra året var väldigt tufft , med allt som hände med mina skador och förändringarna i klubben , men nu har vi en bra känsla .
Truppen är bra och killarna har roligt , träningen är bra .
Förhoppningsvis kan vi gå framåt nu , lägga förra säsongen bakom oss och lyckas bra " .
Kvinnor sover dåligt på grund av rädsla för pensionsbesparingarna
Trots att deltagarna i undersökningen hade en tydlig bild av hur de vill bli omhändertagna var det få som pratade med sina familjemedlemmar om det .
Ungefär hälften av personerna som deltog i den landsomfattande studien sade att de hade pratat med sina makar om kostnaden för långtidsvård .
Bara 10 % sade att de hade talat med sina barn om det .
" Folk vill att en familjemedlem ska ta hand om dem , men de tar inte steget och pratar om det , sade Holly Snyder , vice ordförande för livförsäkringar på Nationwide .
Så här kan du börja .
Tala med din make / maka och barnen : Du kan inte förbereda din familj på att ge dig vård om du inte talar om hur du vill ha det i god tid .
Arbeta med din rådgivare och din familj och diskutera var och hur du vill ha vård . Dina val kan ha stor betydelse för kostnaderna .
Ta hjälp av din ekonomiska rådgivare : Din rådgivare kan också hjälpa dig att hitta ett sätt att betala för kostnaderna .
Dina val av finansiering för långtidsvård kan omfatta en traditionell försäkringslösning för långtidsvård , en hybridlösning med livförsäkring med kontantvärde för att täcka kostnaderna , eller en självförsäkring med egna medel , om du har råd .
Upprätta juridiska handlingar : Undvik juridiska strider från början .
Upprätta en vårdfullmakt , så att du kan utse en betrodd person som ser över din medicinska vård och ser till att vårdpersonalen följer dina önskningar , om du blir oförmögen att kommunicera .
Överväg också en fullmakt för din ekonomi .
Du väljer då en betrodd person som kan fatta ekonomiska beslut i ditt ställe och se till att dina räkningar blir betalda om du själv är oförmögen .
Glöm inte bort detaljerna : Tänk dig att du har en åldrig förälder som hamnar i ett akut medicinskt tillstånd och är på väg till sjukhuset .
Skulle du då kunna svara på frågor om mediciner och allergier ?
Skriv ner sådana detaljer så att du är redo .
" Det är inte bara ekonomin som står på spel , men vilka är läkarna ? " , frågade Martin .
" Vilka mediciner är det ?
Vem tar hand om hunden ?
Se till att ha planen klar " .
Man beskjuten flera gånger med luftgevär i Ilfracombe
En man blev beskjuten flera gånger med luftgevär när han promenerade hem från en utekväll .
Offret , som är i 40 @-@ årsåldern , befann sig i området Oxford Grove i Ilfracombe i Devon när han blev skjuten i bröstet , buken och handen .
Polisen beskriver skjutningen , som ägde rum ca 02 : 30 , som en " enstaka händelse " .
Offret såg inte sin angripare .
Skadorna är inte livshotande , och polisen uppmanar vittnen att höra av sig .
Jordbävningar och tsunamier i Indonesien
Minst 384 människor har dödats i en kraftfull jordbävning och tsunami som drabbade staden Palu i Indonesien i fredags . Det uppger tjänstemän . Dödssiffran förväntas stiga .
Kommunikationerna är utslagna , och räddningspersonal har ännu inte kunnat få någon information från förvaltningsområdet Donggala , ett område norr om Palu som ligger närmare jordbävningens epicentrum . Jordbävningen mätte 7,5 på Richterskalan .
Fler än 16 000 människor evakuerades från Palu efter katastrofen .
Här är några fakta om Palu och Donggala , som ligger på ön Sulawesi :
Palu är huvudort i provinsen Centrala Sulawesi , och ligger i en trång bukt på västkusten av ön Sulawesi . Stadens befolkning uppskattades till 379 800 personer 2017 .
Staden firade sitt 40 @-@ årsjubileum när jordbävningen och tsunamin slog till .
Donggala är ett förvaltningsområde som sträcker sig längs mer än 300 km av nordvästra Sulawesis kust .
Förvaltningsområdet , som är en administrativ region under en provins , hade 2017 en befolkning som uppskattades till 299 200 personer .
Stöttepelarna i provinsen Centrala Sulawesis ekonomi är fiske och jordbruk . Det gäller särskilt kustregionen Donggala .
Nickelgruvdrift är också betydelsefull i provinsen , men den ligger huvudsakligen koncentrerad till Morowali , på motsatta kusten av Sulawesi .
Palu och Donggala har drabbats av tsunamier flera gånger de senaste hundra åren , enligt Indonesiens myndighet för katastrofhantering .
1938 dödades fler än 200 personer av en tsunami som förstörde hundratals hus i Donggala .
Även 1996 drabbades västra Donggala av en tsunami som dödade nio personer .
Indonesien ligger i den cirkumpacifiska seismiska eldringen , som ofta drabbas av jordbävningar .
Här följer några av de största jordbävningarna och tsunamierna under senare år :
2004 : En stor jordbävning vid indonesiska Aceh @-@ provinsens västkust på norra Sumatra den 26 december utlöste en tsunami som drabbade 14 länder . 226 000 människor dog längs Indiska Oceanens kuster . Mer än hälften av dem var i Aceh .
2005 : En rad kraftiga jordbävningar drabbade Sumatras västkust i slutet av mars och början av april .
Hundratals människor dog på ön Nias , utanför Sumatras kust .
2006 : En jordbävning med magnituden 6,8 på Richterskalan slog till söder om Java , Indonesiens folkrikaste ö , och utlöste en tsunami som slog in över den södra kusten och dödade nästan 700 personer .
2009 : En jordbävning med magnituden 7,6 slog till nära staden Padang , huvudort i provinsen Västra Sumatra .
Mer än 1 100 människor dog .
2010 : En jordbävning med magnituden 7,5 slog till mot en av Mentawaiöarna utanför Sumatra . En tsunami på upp till tio meter utlöstes . Dussintals byar förstördes och runt 300 personer dödades .
2016 : En grund jordbävning drabbade förvaltningsområdet Pidie Jaya i Aceh och orsakade förstörelse och panik , då folk påmindes om förödelsen vid den dödliga jordbävningen och tsunamin 2004 .
Den här gången utlöstes ingen tsunami , men mer än 100 personer dödades av byggnader som rasade samman .
2018 : Stora jordbävningar drabbade den indonesiska turistön Lombok . Mer än 500 personer dog , de flesta på den norra sidan av ön .
Jordbävningen förstörde tusentals byggnader , och tusentals turister blev tillfälligt strandsatta .
Sarah Palins äldste son gripen anklagad för våld i hemmet
Track Palin , äldste son till den tidigare Alaskaguvernören och vicepresidentkandidaten Sarah Palin , har gripits anklagad för misshandel .
Palin , som är 29 år och från Wasilla i Alaska , greps misstänkt för våld i hemmet , för att ha lagt sig i en anmälan om våld i hemmet och för att ha motsatt sig gripandet , enligt en rapport som släpptes på lördagen av Alaskas delstatspolis .
Enligt polisrapporten ska han ha tagit telefonen ifrån en kvinnlig bekant som försökte ringa polisen och anmäla de påstådda brotten .
Palin sitter frihetsberövad i Mat @-@ Su @-@ häktet och hålls mot borgen på 500 dollar som ska betalas om den misstänkte bryter mot borgensvillkoren , enligt tv @-@ kanalen KTUU .
Han framträdde i rätten i lördags och förklarade sig " garanterat icke skyldig " när han blev ombedd att uppge sin inställning , enligt tv @-@ kanalen .
Palin misstänks för tre fall av mindre allvarliga brott enligt klass A , vilket innebär att han kan få fängelse i upp till ett år och 250 000 dollar i böter .
Han har också anklagats för ett fall av mindre allvarligt brott enligt klass B , vilket straffas med en dag i fängelse och 2 000 dollar i böter .
Det är inte första gången Palin anklagas för brott .
I december 2017 anklagades han för våld mot sin far , Todd Palin .
Hans mor , Sarah Palin , ringde polisen för att anmäla det påstådda brottet .
Fallet handläggs nu av Alaskas veterandomstol .
I januari 2016 anklagades han för våld i hemmet , för att ha lagt sig i anmälan av våld i hemmet och för innehav av vapen under påverkan i samband med den händelsen .
Hans flickvän anklagar honom för att ha slagit henne i ansiktet .
Sarah Palin fick kritik av veterangrupper 2016 efter att hon hade kopplat sin sons våldsamma beteende till posttraumatiskt stressyndrom , som härrör från hans militärtjänst i Irak .
Jordbävning och tsunami i Indonesien : hundratals döda
Minst 384 människor har dött efter att en jordbävning drabbade ön Sulawesi i Indonesien i fredags .
Jordbävningen , som mätte 7,5 på Richterskalan , utlöste en tsunami och har förstört hundratals hem .
Elförsörjningen och kommunikationerna ligger nere , och dödssiffrorna förväntas stiga de närmaste dagarna .
Jordbävningen slog till strax utanför centrala Sulawesi , som ligger nordost om Indonesiens huvudstad Jakarta .
Filmer som visar när den slog till cirkulerar nu på sociala medier .
Hundratals människor hade samlats till en strandfestival i staden Palu när tsunamin slog in över kusten .
Federala åklagare yrkar på sällsynt dödsstraff för en misstänkt för terrorangrepp i New York
Federala åklagare i New York yrkar på dödsstraff för Sayfullo Saipov , den misstänkte för terrorattentatet i New York som dödade åtta personer . Det är ett sällsynt straff som inte har verkställts för ett federalt brott i delstaten sedan 1953 .
Saipov , 30 , ska ha använt en hyrlastbil från bygg- och inredningskedjan Home Depot för att utföra ett angrepp på en cykelväg längs West Side Highway på nedre Manhattan . Han mejade ner fotgängare och cyklister i sin väg vid attacken , som ägde rum i oktober .
För att motivera en dödsdom måste åklagarna bevisa att Saipov " avsiktligen " dödade de åtta offren och " avsiktligen " orsakade allvarlig kroppsskada , enligt den avsiktsförklaring om dödsstraff som lämnades in i Southern District i New York .
Båda anklagelsepunkterna kan innebära en dödsdom , enligt domstolshandlingen .
Några veckor efter attacken åtalades Saipov av en federal jury på 22 punkter , däribland åtta fall av mord för att stötta beskyddarverksamhet , vilket ofta används av federala åklagare i mål om organiserad brottslighet , samt misshandel och förstörelse av motorfordon .
Attacken krävde " omfattande planering och uppsåt " , sade åklagarna , och beskrev samtidigt sättet som Saipov utförde den på som " avskyvärd , grym och omänsklig " .
Sayfullo Habibullaevic Saipov har orsakat familj och vänner till Diego Enrique Angelini , Nicholas Cleves , Ann @-@ Laure Decadt , Darren Drake , Ariel Erlij , Hernan Ferruchi , Hernan Diego Mendoza och Alejandro Damian Pagnucco skada och förlust " , står det i avsiktsförklaringen .
Fem av offren var turister från Argentina .
New Yorks södra distrikt har inte åtalat i ett mål där det yrkas på dödsstraff på ett decennium .
Den tilltalade , Khalid Barnes , fälldes för mord på två knarklangare , men dömdes slutligen till livstids fängelse i september 2009 .
Senast dödsstraffet verkställdes i ett federalt mål i New York var 1953 . Det gifta paret Julius och Ethel Rosenberg avrättades efter att ha dömts för stämpling till spioneri för Sovjetunionen under det kalla kriget två år tidigare .
Paret Rosenberg avrättades båda i elektriska stolen den 19 juni 1953 .
Saipov , som är uzbekisk medborgare , uppvisade enligt domstolsdokumenten en brist på ånger under de dagar och månader som följde på attacken .
Enligt polisen uppgav han för utredarna att han var nöjd med vad han hade gjort .
Enligt åtalet berättade Saipov för myndigheterna att han fick inspiration till attacken efter att ha tittat på IS @-@ filmer på sin telefon .
Han bad också om att få sätta upp IS @-@ flaggan på sitt sjukhusrum , uppgav polisen .
Han har förklarat sig icke skyldig till de 22 anklagelsepunkterna i åtalet .
David Patton är en av de federala offentliga försvarare som företräder Saipov . Han uppgav att de är " givetvis besvikna " på åklagarsidans beslut .
" Vi anser att beslutet att yrka på dödsstraff i stället för att gå med på livstids fängelse utan möjlighet till villkorlig frigivning om den tilltalade erkänner sig skyldig bara förlänger traumat som dessa händelser har orsakat för samtliga inblandade " , sade Patton .
Saipovs team av försvarare hade tidigare bett åklagarna att inte yrka på dödsstraff .
Parlamentsledamot från Tories säger att NIGEL FARAGE borde få ansvar för Brexitförhandlingarna
Nigel Farage lovade att " mobilisera folkets armé " i dag under en protest på Tories konferens .
Den tidigare UKIP @-@ ledaren sade att politikerna måste " känna hettan " från EU @-@ skeptikerna , när en av Theresa Mays egna parlamentsledamöter föreslog att han skulle leda förhandlingarna med EU .
Den konservative ledamoten Peter Bone sade vid marschen i Birmingham att Storbritannien redan " skulle ha gått ur " om Nigel Farage hade varit Brexitminister .
Men den utmaning som Theresa May står inför när det gäller att få de djupt delade anhängarna att försonas har förvärrats av EU @-@ positiva torymedlemmar , som har anslutit sig till en separat protest mot Brexit i staden .
Premiärministern kämpar för att hålla sin kompromissplan , Chequers @-@ avtalet , vid liv under angrepp från Brexitanhängare , personer som vill stanna i unionen och EU självt .
Hennes allierade har insisterat på att hon bör trycka på och försöka få till ett avtal med Bryssel trots bakslaget , och tvinga EU @-@ skeptiker och Labourpartiet att välja mellan hennes paketlösning och " kaos " .
Bone sade vid ett massmöte som hade organiserats av organisationen Leave Means Leave i Solihull att han ville " spola Chequers @-@ avtalet " .
Han antydde att Nigel Farage borde ha gjorts till jämlike och fått ansvarsområden vid förhandlingarna med Bryssel .
" Om han hade stått vid rodret så hade vi varit ute vid det här laget " , sade han .
Peter Bone , som representerar distriktet Wellingborough i parlamentet , tillade : " Jag kommer att stå upp för Brexit , men vi måste spola Chequers @-@ avtalet " .
Han tydliggjorde sitt motstånd mot EU och sa : " Vi har inte utkämpat världskrig för att bli undersåtar .
Vi vill stifta våra egna lagar i vårt eget land " .
Bone avfärdade påståendena om att den allmänna opinionen skulle ha förändrats sedan folkomröstningen 2016 : " Tanken att britterna skulle ha ändrat sig och nu vill stanna kvar är helt osann " .
Brexitanhängaren Andrea Jenkyns från Torypartiet var också med på marschen och talade med journalisterna . " Jag vill bara säga : " Premiärministern , lyssna till folket " .
Chequers @-@ avtalet är impopulärt hos allmänheten , oppositionen kommer inte att rösta för det , det är impopulärt i partiet och hos våra valarbetare som är ute på gatorna och ser till att vi blir valda .
Lägg undan Chequers @-@ avtalet och börja lyssna " .
Och hon tillade ett skarpt budskap riktat till Theresa May : " Premiärministrar får behålla sina jobb när de håller sina löften " .
Nigel Farage sade vid mötet att politikerna måste få " känna hettan " om de skulle svika beslutet som fattades i och med folkomröstningen 2016 .
" Nu handlar det om förtroendet mellan oss , det vill säga folket , och den politiska klassen " , sade han .
" De försöker svika Brexit , och vi är här i dag för att säga till dem : " Vi tänker inte låta er komma undan med det " . "
Inför den entusiastiska folkmassan tillade han : " Jag vill att ni ska få vår politiska klass , som är nära att svika Brexit , att känna hettan .
Vi mobiliserar folkets armé i det här landet som gav oss seger i Brexit , och vi kommer inte att vila förrän vi har blivit ett självständigt , självstyrande och stolt Storbritannien " .
Samtidigt marscherade EU @-@ anhängare genom Birmingham och höll sedan ett två timmar långt massmöte i centrala staden .
En grupp aktivister viftade med baner med texten " Torymedlemmar mot Brexit " efter att gruppen lanserades i helgen .
Labourparlamentarikern Lord Adonis från Överhuset hånade de konservativa för säkerhetsproblemen de stötte på med en partiapp när konferensen öppnade .
" Det är de här människorna som säger att de kan ha IT @-@ system på plats och all teknik för Kanada plus plus plus @-@ avtalet , för friktionslösa gränser och frihandel utan gränser i Irland " , tillade han .
" Det är en ren fars .
Det finns ingen god Brexit " , tillade han .
Warren planerar en " ordentlig funderare " om att kandidera till presidentposten
Den amerikanska senatorn Elizabeth Warren säger att hon ska ta sig en " ordentlig funderare om att kandidera till presidentposten " efter valen i november .
Tidningen Boston Globe rapporterar att demokraten från Massachusetts talade om sin framtid under ett stadshusmöte i västra Massachusetts i lördags .
Warren har ofta kritiserat president Donald Trump , och ställer nu upp för omval i november mot den republikanske delstatsrepresentanten Geoff Diehl , som var biträdande ordförande i Donald Trumps kampanj i Massachusetts 2016 .
Hon har varit föremål för spekulationer om att hon kanske tar sig an Donald Trump 2020 .
Evenemanget på lördag eftermiddag i Holyoke var hennes 36:e stadshusmöte med väljarna sedan Donald Trump tillträdde .
En person frågade henne om hon planerade att kandidera till presidentposten .
Warren svarade att det är dags " för kvinnor att åka till Washington för att reparera vår trasiga regering . Det innebär en kvinna på toppen " .
En person gripen för dödsskjutningen av basketspelaren Sims från LSU
Polisen i Baton Rouge i Louisiana tillkännagav på lördagen att en misstänkt hade gripits för dödsskjutningen av LSU @-@ basketspelaren Wayde Sims på fredagen .
Polisen i Baton Rouge tillkännagav att Dyteon Simpson , 20 , hade gripits vid en presskonferens klockan 11 : 00 för ET .
De hade släppt en film av skjutningen på fredagen för att få hjälp att identifiera en man som syns på bilderna .
20 @-@ årige Sims sköts till döds nära Southern Universitys campus tidigt på fredagen .
" Wayde Sims blev skottskadad i huvudet och dog slutligen av detta " , berättade polischefen Murphy J. Paul för medierna på lördagen via nyhetssajten 247 sports .
Wayde gick emellan för att försvara sin vän och blev skjuten av Simpson .
Simpson förhördes och erkände att han hade varit på platsen och haft ett vapen , och han erkände att han hade skjutit Wayde Sims .
Simpson greps utan några incidenter och fördes till häktet vid polisen i East Baton Rouge .
Sims var juniorspelare , 198 cm lång och växte upp i Baton Rouge . Han spelade i 32 matcher med 10 starter förra säsongen , och snittade på 17,4 minuter , 5,6 poäng och 2,9 returer per match .
Rysslands Grand Prix : Lewis Hamilton närmar sig världsmästartiteln efter det att teamorder gav honom vinst över Sebastian Vettel
Från det ögonblick då Valtteri Bottas kvalificerade sig före Lewis Hamilton på lördagen stod det klart att Mercedes " teamorder skulle spela en stor roll i loppet .
Bottas fick en bra start och hängde nästan ut Hamilton på tork när han försvarade sin position under de första två varven , och bjöd in Vettel att angripa sin lagkamrat .
Vettel gick i depå först och lät Hamilton köra in längst bak i klungan , vilket bör ha varit avgörande .
Mercedesen gick i depå ett varv senare och kom ut bakom Vettel , men Hamilton gick framåt efter lite hjul @-@ mot @-@ hjul @-@ action där Ferrari @-@ föraren motvilligt lämnade insidan fri med risk för att bjuda på plats efter ett dubbeldrag för att försvara sig i det tredje kurvan .
Max Verstappen startade i den bakre raden och låg sjua i slutet av första varvet på sin 21 @-@ årsdag .
Han ledde sedan en stor del av loppet och höll i däcken för att nå en snabb målgång och köra om Kimi Raikkonen och bli fyra .
Till slut kom han i depån på 44:e varvet men lyckades inte höja tempot under de kvarvarande åtta varven när Raikkonen gick upp på fjärde plats .
Det är en svår dag , eftersom Valtteri gjorde ett fantastiskt jobb hela helgen och var en riktig gentleman som släppte förbi mig .
Teamet har gjort ett exceptionellt jobb och fått en etta och en tvåa " , sade Hamilton .
Riktigt dåligt kroppsspråk
President Donald Trump hånade senator Dianne Feinstein vid ett massmöte på lördagen , för att hon vidhåller att hon inte har läckt brevet från Christine Blasey Ford i vilket Brett Kavanaugh , som är nominerad till domare i Högsta Domstolen , anklagas för sexuella övergrepp .
Presidenten , som talade vid ett massmöte i West Virginia , tog inte direkt upp vittnesmålet från Ford inför senatens justitieutskott . I stället kommenterade han att det som pågick i senaten visade att folk var " elaka , otäcka och lögnaktiga " .
" Det enda som kunde hända och det fina som har hänt de senaste dagarna i senaten , när man ser ilskan , när man ser folk som är arga , elaka , otäcka och lögnaktiga " , sade han .
" Man ser pressmeddelanden och läckor och så säger de : " Nej , jag har inte gjort det .
Jag har inte gjort det " .
Kommer ni ihåg ?
Har du läckt , Dianne Feinstein ?
Kommer ni ihåg hennes svar ? " Har du läckt dokumentet ? " " Åh , vadå ? "
Åh , nej .
Jag har inte läckt det " .
Vänta lite nu .
" Har vi läckt ... Nej , vi har inte läckt något " " , tillade han , och imiterade senatorn .
Brevet med detaljer om Fords anklagelser mot Kavanaugh skickades till Feinstein i juli , och läcktes i september , men Feinstein förnekade att läckan skulle ha kommit från hennes kontor .
" Jag har inte mörkat Fords anklagelser , jag har inte läckt hennes berättelse " , sade Feinstein till kommittén enligt tidningen The Hill .
" Hon bad mig att hålla detta konfidentiellt , och jag höll det konfidentiellt , som hon önskade " .
Men hennes dementi verkar inte ha passat presidenten , som under lördagskvällens möte kommenterade det så här : " Jag ska säga er en sak . Det där var verkligen dåligt kroppsspråk .
Hon kanske inte har gjort det , men det där var det sämsta kroppsspråket jag har sett " .
Presidenten fortsätter att stötta kandidaten till Högsta Domstolen , som har blivit anklagad för sexualbrott av tre kvinnor , och han antydde att demokraterna använde anklagelserna för sina egna syften .
" De är fast beslutna att ta tillbaka makten med alla nödvändiga medel .
Man ser deras elakhet och vidrighet . De bryr sig inte om vem de skadar , vem de måste köra över för att få makt och kontroll " , sade presidenten enligt den digitala nyhetssajten Mediaite .
Elite League : Dundee Stars @-@ Belfast Giants 5 @-@ 3
Patrick Dwyer gjorde två mål för Belfast Giants mot Dundee
Dundee Stars sonade fredagens förlust i Elite League mot Belfast Giants genom att vinna returmatchen med 5 @-@ 3 i Dundee på lördagen .
Belfast Giants fick en tidig tvåmålsledning genom Patrick Dwyer och Francis Beauvillier .
Mike Sullivan och Jordan Cownie kvitterade för hemmalaget innan Dwyer återupprättade Belfast Giants ledning .
Francois Bouchard kvitterade för Dundee innan två mål från Lukas Lundvald Nielsen säkrade segern .
Det var den tredje förlusten i Elite League för säsongen för Adam Keefes lag , som kom bakifrån och slog Dundee med 2 @-@ 1 i Belfast på fredagskvällen .
Det var det fjärde mötet för säsongen för de två lagen , och Belfast Giants hade vunnit de tre tidigare matcherna .
Dwyers öppningsmål kom i den fjärde minuten vid 3 : 35 på assist från Kendall McFaull , och David Rutherford gav assist när Beauvillier fördubblade ledningen fyra minuter senare .
I den intensiva första perioden förde Sullivan hemmalaget tillbaka in i matchen vid 13 : 10 innan Matt Marquardt levererade till Cownie som kvitterade vid 15 : 16 .
Dwyer såg till att Belfast Giants låg i ledningen vid den första pausen när han gjorde sitt andra mål för kvällen i slutet av den första perioden .
Hemmalaget omgrupperade sig och Bouchard kvitterade än en gång med ett mål i power play vid 27 : 37 .
Cownie och Charles Corcoran samarbetade för att hjälpa Nielsen ge Dundee ledningen för första gången i matchen i slutet av andra perioden , och han säkrade vinsten med sitt lags femte halvvägs igenom slutperioden .
Belfast Giants , som nu har förlorat fyra av sina fem senaste matcher , ska spela hemma mot Milton Keynes vid sin nästa match på fredag .
Flygledare dog för att hundratals människor på ett plan skulle kunna fly från jordbävning
En flygledare i Indonesien hyllas nu som en hjälte efter det att han avled när han såg till att ett plan med hundratals människor ombord kunde lyfta säkert .
Mer än 800 personer har dött och många saknas efter det att en stor jordbävning drabbade ön Sulawesi på fredagen och utlöste en tsunami .
Kraftiga efterskalv fortsätter att plåga området och många är fast i bråten i staden Palu .
Men trots att hans kollegor flydde för sina liv vägrade 21 @-@ årige Anthonius Gunawan Agung lämna sin post i det vilt svajande kontrolltornet på flygplatsen Mutiara Sis Al Jufri i Palu .
Han stannade kvar för att se till att Batik Airs flight 6321 , som då befann sig på startbanan , kunde lyfta säkert .
Sedan hoppade han från kontrolltornet när han trodde att det skulle rasa .
Han avled senare på sjukhus .
Talespersonen för Air Navigation Indonesia , Yohannes Sirait , sade att beslutet kan ha räddat hundratals människors liv , enligt den australiska tv @-@ kanalen ABC News .
" Vi ordnade med en helikopter från Balikpapan på Kalimantan för att ta honom till ett större sjukhus i en annan stad .
Tyvärr avled han i morse innan helikoptern kom fram till Palu .
Vi är förkrossade över att få höra detta " , tillade han .
Samtidigt befarar myndigheterna att dödssiffran kan stiga till över tusen personer . Landets katastrofhjälpsmyndighet säger att det är begränsad åtkomst till städerna Donggala , Sigi och Boutong .
" Dödssiffran tros fortsätta öka eftersom det fortfarande är många kroppar kvar i ruinerna , och många har inte kunnat nås " , sade Sutopo Purwo Nugroho , en talesperson för myndigheten .
Upp till sex meter höga vågor har ödelagt Palu , där en massbegravning kommer att hållas på söndag .
Militära och kommersiella flygplan flyger in hjälp och förnödenheter .
Den 35 @-@ åriga mamman Risa Kusuma sade till Sky News : " Varje minut kommer en ambulans med döda kroppar .
Det är ont om rent vatten .
Minimarknaderna plundras överallt " .
Jan Gelfand , chef för Internationella Röda Korset i Indonesien , sade till CNN : " Det indonesiska Röda Korset kämpar för att hjälpa överlevande , men vi vet inte vad de kommer att mötas av där .
Detta är redan en tragedi , men det kan bli mycket värre " .
Indonesiens president Joko Widodo anlände till Palu på söndagen och sade till landets militär : " Jag ber er alla att arbeta dag och natt för att slutföra alla uppgifter som är relaterade till evakueringen .
Är ni redo ? " enligt CNN .
Indonesien drabbades tidigare i år av jordbävningar på Lombok , där mer än 550 personer omkom .
Flygplanskrasch i Mikronesien : Air Niugini uppger nu att en man saknas efter att ett flygplan störtat i en lagun
Flygbolaget som ansvarar för det plan som störtade i en lagun i Mikronesien i Stilla Havet uppger nu att en man saknas . Tidigare sades det att alla 47 passagerare och besättningen hade utrymts från det sjunkande planet och befann sig i säkerhet .
Air Niugini sade i ett pressmeddelande att en manlig passagerare fortfarande saknades på lördagseftermiddagen .
Flygbolaget sade att det arbetade tillsammans med lokala myndigheter , sjukhus och utredare för att försöka hitta mannen .
Flygbolaget svarade inte genast på frågorna om fler detaljer om passageraren , som exempelvis hans ålder och nationalitet .
Lokala båtar hjälpte till att rädda de andra passagerarna och besättningen efter det att planet störtade i vattnet då det försökte landa på flygplatsen på Chuuköarna .
Tjänstemän uppgav på fredagen att sju personer hade förts till sjukhus .
Flygbolaget uppgav att sex passagerare var kvar på sjukhuset på lördagen och att deras tillstånd var stabilt .
Det är ännu oklart vad som orsakade kraschen och hur händelseförloppet såg ut .
Flygbolaget och den amerikanska flottan uppgav båda att planet landade i lagunen utan att nå landningsbanan .
Vissa vittnen trodde att planet gled förbi landningsbanan .
Den amerikanske passageraren Bill Jaynes sade att planet flög in mycket lågt .
" Det är extremt bra " , sade Jaynes .
Jaynes sade att han och andra lyckades vada genom midjedjupt vatten till nödutgångarna på det sjunkande planet .
Han sade att kabinpersonalen fick panik och skrek , och att han fick en mindre skallskada .
Den amerikanska flottan sade att sjömän som arbetade i närheten med att utveckla ett skeppsvarv också hjälpte till i räddningsarbetet genom att använda en uppblåsbar båt för att köra folk i land innan planet sjönk i det 30 meter djupa vattnet .
Data från Aviation Safety Network visar att 111 personer har omkommit i olyckor med flygbolag som är registrerade i Papua Nya Guinea de senaste två åren , men Air Niugini har inte varit inblandat i någon av dem .
Analytiker ritar upp en tidslinje för natten då en kvinna brändes levande
Åklagarsidan avslutade på lördagen sin plädering i den andra rättegången mot en man som anklagas för att ha bränt en kvinna i Mississippi levande 2014 .
Det amerikanska justitiedepartementets analytiker Paul Rowlett talade i timmar som expertvittne på området underrättelseanalys .
Han förklarade för juryn hur han hade använt mobiltelefonlistor för att pussla ihop den 29 @-@ årige tilltalade Quinton Tellis och det 19 @-@ åriga offret Jessica Chambers rörelser den natten hon dog .
Rowlett sade att han hade fått lokaliseringsuppgifter från flera mobiltelefoner som visade att Tellis var med Chambers den kvällen hon dog , vilket motsäger hans tidigare påståenden , rapporterade nyhetstidningen The Clarion Ledger .
När uppgifterna visade att hans mobiltelefon var tillsammans med Chambers mobiltelefon under den tidsperiod han sade att han hade varit med sin vän Michael Sanford , så gick polisen för att tala med Sanford .
Sanford vittnade i lördags och sade att han inte var i staden den dagen .
När åklagarna frågade om Tellis sade sanningen när han sade att han var i Sanfords lastbil den kvällen , så sade Sanford att han " ljuger , för min lastbil var i Nashville " .
En annan motsägelse var att Tellis uppgav att han hade känt Chambers i ungefär två veckor när hon dog .
Mobiltelefonlistor visade att de bara hade känt varandra i en vecka .
Rowlett sade att Tellis en tid efter Chambers " död raderade Chambers " textmeddelanden , samtal och kontaktinformation från sin telefon .
" Han suddade ut henne från sitt liv " , sade Hale .
Försvaret planeras påbörja sitt slutanförande på söndag .
Domaren sade att han väntade sig att prövningen skulle överlämnas till juryn senare samma dag .
The High Breed : Vad är medveten hiphop ?
En hiphop @-@ trio vill utmana den negativa bilden av genren genom att fylla sin musik med positiva budskap .
The High Breed från Bristol tycker att hiphopen har kommit långt bort från sitt ursprung i politiska budskap och att angripa sociala frågor .
De vill gå tillbaka till rötterna och göra medveten hiphop populär igen .
Artister som The Fugees och Common har nyligen fått ett uppsving i Storbritannien genom artister som Akala och Lowkey .
En svart igen ? !
En barnflicka i New York stämmer ett par på grund av uppsägning efter ett " rasistiskt " textmeddelande
En barnflicka i New York stämmer ett par för diskriminerande uppsägning efter att hon fått ett felskickat textmeddelande från modern , som klagade över att hon var " en svart igen " .
Paret förnekar att de skulle vara rasister och jämför stämningen med " utpressning " .
Tvåbarnsmamman Lynsey Plasco @-@ Flaxman uttryckte förskräckelse när hon förstod att den nya barnflickan Giselle Maurice var svart , då hon kom till sin första arbetsdag 2016 .
" NEEEEEEEEEEEJ INTE EN SVART IGEN " , skrev Lynsey Plasco @-@ Flaxman i ett sms till sin man .
Men i stället för att skicka det till sin man skickade hon det till Giselle Maurice , två gånger .
Efter att hon hade insett sitt misstag var Plasco @-@ Flaxman " illa till mods " , och gav Maurice sparken , och hävdade att deras tidigare barnflicka , som var afroamerikan , hade gjort ett dåligt jobb och att hon i stället förväntade sig en filippinsk kvinna , enligt New York Post .
Maurice fick betalt för en dags arbete och skickades hem i taxi .
Nu stämmer hon paret för att få kompensation för avskedandet . Hon begär ersättning i storleksordningen 350 dollar per dag för jobbet hon från början anställdes för att göra , som skulle vara i sex månader och där hon skulle bo hos paret . Dock hade hon inget kontrakt .
" Jag vill visa dem att man inte gör så " , sade hon till New York Post på fredagen . " Jag vet att det är diskriminering " .
Paret slår ifrån sig anklagelserna om att de skulle vara rasister och säger att det enda raka var att avsluta Giselle Maurices anställning . De var oroliga för att de inte skulle kunna lita på henne när de hade förolämpat henne .
" Min fru hade skickat henne något som hon inte menade .
Hon är inte rasist .
Vi är inte rasister " , sade maken Joel Plasco till New York Post .
" Men skulle du anförtro dina barn till någon som du hade varit oförskämd mot , även om det var av misstag ?
Din nyfödda bebis ?
Allvarligt talat " .
Plasco jämförde stämningen med " utpressning " och sade att hans fru skulle föda barn två månader senare och befann sig i en " mycket svår situation " .
" Ska man ge sig på en sådan person ?
Det är inte särskilt trevligt gjort " , tillade investeringsbankiren Plasco .
Rättsprocessen pågår fortfarande , men den allmänna opinionen har snabbt fördömt paret på sociala medier och kritiserar dem för deras beteende och resonemang .
Paddington @-@ förläggarna trodde inte att läsarna skulle kunna relatera till en talande björn , avslöjar ett nytt brev
Paddington @-@ författaren Michael Bonds dotter Karen Jankel , som föddes strax efter det att boken blev antagen , kommenterade brevet så här : " Det är svårt att tänka sig in i hur det var för en person som läste den för första gången innan den gavs ut .
Det är väldigt roligt , med tanke på det vi nu vet om Paddingtons stora framgång " .
Hon berättade att hennes pappa , som hade arbetat som kameraman på BBC innan han fick inspiration av en liten leksaksbjörn att skriva barnboken , hade varit optimistisk när hans arbete förkastades . Hon tillade att 60 @-@ årsjubiléet av den första utgåvan var " bitterljuvt " efter hans död förra året .
Hon beskriver att Paddington var en " mycket viktig medlem av vår familj " , och tillade att hennes far var stolt i det tysta över sin slutliga framgång .
" Han var ganska tystlåten av sig , och inte någon skrytsam person " , sade hon .
" Men Paddington var så verklig för honom , det var nästan som att ha ett barn som lyckas med något . Man blir stolt över barnet även om det inte är man själv som har åstadkommit det .
Jag tror att han såg Paddingtons framgångar lite på det sättet .
Även om det var hans skapelse och hans fantasi brukade han alltid ge Paddington själv äran " .
Min dotter skulle dö , och jag fick ta farväl i telefonen
När hon landade hade hennes dotter förts i ilfart till sjukhuset Louis Pasteur 2 i Nice , där läkarna arbetade förgäves för att rädda hennes liv .
" Nad ringde regelbundet för att säga att det var riktigt illa , och att man inte väntade sig att hon skulle klara sig " , sade mrs Ednan @-@ Laperouse .
" Sedan fick jag ett samtal från Nad som sade att hon skulle dö inom två minuter och att jag måste ta farväl av henne .
Och det gjorde jag .
Jag sa : " Jag älskar dig så mycket , Tashi , min älskling .
Jag kommer till dig snart .
Jag kommer till dig .
Medicinerna som läkarna hade gett henne för att hålla hennes hjärta vid liv ebbade långsamt ut och lämnade hennes kropp .
Hon hade dött strax innan och nu släcktes allting ned .
Jag fick bara sitta där och vänta och veta att allt detta hände .
Jag kunde inte tjuta eller skrika eller gråta , eftersom jag var omgiven av familjer och människor .
Jag var tvungen att ta mig samman " .
Slutligen gick mrs Ednan @-@ Laperouse , som nu sörjde förlusten av sin dotter , ombord på planet tillsammans med de andra passagerarna , som var helt omedvetna om den svåra prövning hon gick igenom .
" Ingen visste om det " , sade hon .
" Jag böjde ned huvudet , och tårarna rann hela tiden .
Det är svårt att förklara , men på flyget kände jag en överväldigande medkänsla för Nad .
Att han behövde min kärlek och min förståelse .
Jag visste hur mycket han älskade henne " .
Sörjande kvinnor sätter upp vykort för att förebygga självmord på bro
Två kvinnor som har förlorat närstående på grund av självmord arbetar för att förhindra att andra tar sina liv .
Sharon Davis och Kelly Humphreys har satt upp kort på en bro i Wales med inspirerande budskap och telefonnummer som man kan ringa för att få stöd .
Sharon Davis ' son Tyler var 13 år när han började lida av depression , och tog sitt liv när han var 18 .
" Jag vill inte att någon förälder ska behöva må så dåligt som jag gör varje dag " , säger hon .
Sharon Davis är 45 år och bor i Lydney . Hon berättar att hennes son var en lovande kock som hade ett smittande leende .
" Alla visste vem han var på grund av hans leende .
De sade att hans leende lyste upp rummet " .
Men han slutade arbeta innan han dog , eftersom han befann sig " på en väldigt mörk plats " .
Tylers bror , som då var 11 år , var den som hittade sitt syskon när han hade tagit livet av sig 2014 .
Sharon Davis säger : " Jag oroar mig hela tiden för följdverkningar " .
Sharon Davis skapade korten " för att människor ska veta att det finns folk man kan gå och prata med , även om det är en vän .
Sitt inte tyst , prata om det " .
Kelly Humphreys , som har varit vän med Sharon Davies i åratal , miste sin partner sedan 15 år , Mark , en tid efter hans mammas död .
" Han hade inte sagt att han kände sig nedstämd eller deprimerad eller någonting " , säger hon .
" Några dagar innan jul märkte vi att han betedde sig annorlunda .
På juldagen befann han sig på botten . När barnen öppnade sina julklappar hade han inte ögonkontakt med dem eller nåt " .
Hon säger att hans död var ett mycket hårt slag för dem , men de måste ta sig igenom det . " Det river upp ett sår i familjen .
Det sliter sönder oss .
Men vi måste kämpa vidare allihop " .
Om du också har det svårt kan du ringa organisationen Samaritans gratis på 116 123 ( Storbritannien och Irland ) , e @-@ posta till jo @ samaritans.org eller gå in på Samaritans hemsida här .
Brett Kavanaughs framtid står på spel när FBI inleder utredning
" Jag tänkte att om vi kunde åstadkomma något som liknar det han bad om - en utredning som är begränsad i tid och omfattning - så kunde vi kanske få lite enighet " , sade Jeff Flake på lördagen . Han tillade att han fruktade att kommittén skulle " splittras " på grund av djupt rotade partsskiljaktigheter .
Varför ville inte Kavanaugh och hans republikanska anhängare att FBI skulle utreda fallet ?
Deras motsträvighet beror helt på tidpunkten .
Mellanårsvalen ska äga rum om bara fem veckor , den 6 november . Om republikanerna gör ett dåligt val , vilket är väntat , kommer de att vara kraftigt försvagade i sina försök att få den man de vill ha vald till landets högsta domstol .
George W. Bush har tagit telefonen och ringt till senatorer för att påverka dem att stötta Kavanaugh , som arbetade åt Bush i Vita huset och genom honom träffade sin fru Ashley , som var personlig sekreterare åt George W. Bush .
Vad händer efter det att FBI lägger fram sin rapport ?
Det blir en omröstning i senaten , där det nu sitter 51 republikaner och 49 demokrater .
Det är fortfarande oklart om Kavanaugh kan få minst 50 röster i senaten , vilket skulle göra att vicepresidenten Mike Pence kan bryta dödläget och bekräfta hans inval i Högsta Domstolen .
Antalet nordkoreanska avhoppare " sjunker " under Kim
Antalet nordkoreaner som hoppar av till Sydkorea har sjunkit sedan Kim Jong @-@ un kom till makten för sju år sedan , säger en sydkoreansk lagstiftare .
Park Byeong @-@ seug , som citerar uppgifter från Sydkoreas återföreningsministerium , säger att 1 127 personer hoppade av förra året , jämfört med 2 706 år 2011 .
Park säger att hårdare gränskontroller mellan Nordkorea och Kina samt högre avgifter till människosmugglare är viktiga orsaker .
Pyongyang har inte kommit med några offentliga kommentarer .
De allra flesta avhoppare från Nordkorea erbjuds slutligen sydkoreanskt medborgarskap .
Enligt Seoul ska mer än 30 000 nordkoreaner ha korsat gränsen illegalt sedan Koreakrigets slut 1953 .
De flesta flyr via Kina , som har längst gräns mot Nordkorea och vars gräns är enklare att korsa än den hårt bevakade demilitariserade zonen ( DMZ ) mellan de båda Koreastaterna .
Kina ser avhopparna som illegala migranter snarare än som flyktingar och skickar ofta tillbaka dem med våld .
Relationen mellan Nord och Syd , som tekniskt sett fortfarande ligger i krig med varandra , har förbättrats markant de senaste månaderna .
Tidigare i månaden träffades ledarna för de två länderna i Pyongyang för samtal med fokus på de fastkörda förhandlingarna om kärnvapennedrustning .
Detta hände efter det historiska mötet i juni mellan USA:s president Donald Trump och Kim Jong @-@ un i Singapore , där de kom överens i generella termer att arbeta för att den koreanska halvön ska bli fri från kärnvapen .
Men på lördagen anklagade Nordkoreas utrikesminister , Ri Yong @-@ ho , de amerikanska sanktionerna för bristen på framgång sedan dess .
" Utan förtroende för USA finns ingen tillit till vår nationella säkerhet , och under sådana omständigheter kan vi absolut inte avväpna oss själva unilateralt först " , sade Ri vid ett tal i FN:s generalförsamling i New York .
Nancy Pelosi kallar Brett Kavanaugh för " hysterisk " , och säger att han är olämplig att tjänstgöra i Högsta Domstolen
Minoritetsledaren i kammaren , Nancy Pelosi , kallade kandidaten till Högsta Domstolen Brett Kavanaugh " hysterisk " och sade att han var temperamentsmässigt olämplig att tjänstgöra i Högsta Domstolen .
Pelosis kommentarer kom i en intervju på lördagen vid Texas Tribune Festival i Austin i Texas .
" Jag kunde inte hjälpa att jag tänkte att om en kvinna hade betett sig så , så skulle hon kallas " hysterisk " " , sade Pelosi om sin reaktion på Kavanaughs vittnesmål inför senatens justitieutskott på torsdagen .
Kavanaugh blev känslomässig när han förnekade anklagelserna om att ha ofredat dr Christine Blasey Ford sexuellt när de båda var tonåringar .
Under sitt öppningsanförande blev Kavanaugh väldigt känslomässigt berörd , och då och då skrek han nästan och rösten stockade sig när han talade om sin familj och sina år i high school .
Han fördömde också uttryckligen demokraterna i kommittén , och sade att anklagelserna mot honom var ett " groteskt och samordnat karaktärsmord " som var organiserat av liberaler som var arga för att Hillary Clinton förlorade presidentvalet 2016 .
Pelosi sade att hon ansåg att Kavanaughs vittnesmål bevisade att han inte kunde tjänstgöra i Högsta domstolen , eftersom det visade att han är partisk till demokraternas nackdel .
" Jag tycker att han diskvalificerar sig själv med sina uttalanden och sättet på vilket han attackerade paret Clinton och demokraterna " , sade hon .
Pelosi tvekade när hon fick frågan om hon skulle försöka ställa Kavanaugh inför riksrätt om han blir invald , och om demokraterna får majoritet i Representanthuset .
" Jag kan säga så här - om han inte säger sanningen till Kongressen eller FBI , då är han inte bara olämplig att sitta i Högsta domstolen , utan också att arbeta i den domstol han är på nu " , sade Pelosi .
Kavanaugh är för närvarande domare i appellationsdomstolen i Washington D.C.
Pelosi tillade att hon som demokrat var orolig för vilka beslut Kavanaugh kan komma att fatta mot sjukvårdsförsäkringslagen Affordable Care Act eller abortmålet Roe vs. Wade , eftersom han anses vara en konservativ domare .
I sina bekräftelseutfrågningar undvek Kavanaugh frågor om huruvida han skulle ändra på vissa beslut av Högsta domstolen .
Det är inte läge för en hysterisk och partisk person att sätta sig i rätten och förvänta sig att vi alla applåderar " , sade Pelosi .
Kvinnor måste stå ut .
Det är en rättfärdig kritik , månader och år av ilska som kokar över , och hon kan inte få ut det utan att gråta .
" Vi gråter när vi blir arga " , sade ms . Steinem till mig 45 år senare .
" Jag tror inte att det är ovanligt . Tror du ? "
Och hon fortsatte : " Jag fick god hjälp av en kvinna som var VD någonstans . Hon sade att hon också grät när hon blev arg , men hade utvecklat en teknik som innebar att när hon blev arg och började gråta sade hon till personen hon talade med : " Du kanske tror att jag är ledsen eftersom jag gråter .
Jag är arg " .
Och så fortsatte hon .
Jag tyckte att det var lysande " .
Tårar är tillåtna för att få utlopp för vrede delvis för att de ofta missförstås i grunden .
Ett av mina tydligaste minnen från ett av mina första jobb på ett mansdominerat kontor , där jag en gång grät av obeskrivlig ilska , var att jag togs i kragen av en äldre kvinna . Det var en kylig chef som jag alltid hade varit lite rädd för , och hon drog mig in i ett trapphus .
" Låt dem aldrig se att du gråter " , sade hon till mig .
" De vet inte att du är rasande .
De tror att du är ledsen och blir glada för att de lyckades trycka till dig " .
Patricia Schroeder , som då var demokratisk kongressledamot från Colorado , hade arbetat med Gary Hart i hans presidentvalskampanjer .
1987 , när Hart ertappades med en utomäktenskaplig affär på en båt som hette Monkey Business och drog sig ur kampanjen , ansåg en mycket frustrerad Schroeder att det inte fanns någon anledning att inte undersöka tanken på att själv ställa upp i presidentvalet .
" Det var inte ett väl genomtänkt beslut " , sade hon med ett skratt till mig 30 år senare .
" Det fanns redan sju andra kandidater . Det sista de behövde var en till .
Någon kallade det för " Snövit och de sju dvärgarna " " .
Eftersom hon var sent ute låg hon efter med pengainsamlingen , och gav löftet att inte gå in som kandidat om hon inte fick ihop 2 miljoner dollar .
Det var ett projekt dömt att misslyckas .
Hon upptäckte att vissa av hennes supportrar som gav 1 000 dollar till män bara gav henne 250 dollar .
" Tror de att jag får rabatt ? " undrade hon .
När hon i ett tal tillkännagav att hon inte skulle inleda en formell presidentvalskampanj blev hon så överväldigad av känslor , tacksamhet mot dem som hade stöttat henne , frustration över systemet som gjorde det så svårt att samla in pengar och rikta sig mot väljare snarare än delegater , och ilska mot sexismen , att rösten stockade sig .
" Man kunde ha trott att jag hade fått ett nervöst sammanbrott " , minns Schröder apropå pressens reaktioner .
" Man kunde ha trott att Kleenex var min företagssponsor .
Jag minns att jag tänkte : " Vad ska de skriva på min gravsten ? "
" Hon grät ? " "
Varför handelskriget mellan USA och Kina kan vara bra för Peking
Öppningstiraden i handelskriget mellan USA och Kina var öronbedövande . Kriget är långt ifrån över , men sprickan mellan länderna kan gynna den kinesiska regeringen på lång sikt , enligt experter .
USA:s president Donald Trump avfyrade det första varningsskottet tidigare i år genom att belägga viktiga kinesiska exportvaror som solpaneler , stål och aluminium med tullar .
Den mest betydelsefulla upptrappningen kom i veckan , med nya tullar på varor för 200 miljarder dollar . Det innebär i praktiken att hälften av allt gods som kommer in i USA från Kina är tullbelagt .
Peking har varje gång svarat med samma mynt . Nyligen slängde man på avgifter på mellan fem och tio procent på amerikanska varor för 60 miljarder dollar .
Kina har lovat att matcha USA:s åtgärder . Världens näst största ekonomi kommer troligen inte att trappa ner inom överskådlig tid .
Att få Washington att backa innebär att böja sig för krav , men att offentligt krypa för USA skulle vara alldeles för genant för Kinas president Xi Jinping .
Experter menar dock att om Peking spelar sina kort rätt kan pressen från USA:s handelskrig ge ett positivt stöd till Kina på lång sikt , genom att minska de två ekonomiernas ömsesidiga beroende av varandra .
" Ett snabbt politiskt beslut i antingen Washington eller Peking kan skapa förutsättningar för ekonomisk panik i endera landet , och det är faktiskt betydligt farligare än betraktarna tidigare har velat erkänna " , säger Abigail Grace , forskningsassistent med fokus på Asien vid tankesmedjan Center for New American Security .
Syrien " redo " för hemvändande flyktingar , enligt utrikesministern
Syrien säger att landet är redo att ta emot frivilligt återvändande flyktingar och vädjar om hjälp för att bygga upp landet , som ligger i ruiner efter det mer än sju år långa kriget .
I ett tal inför FN:s generalförsamling sade utrikesministern Walid al @-@ Moualem att villkoren i landet nu förbättras .
" Situationen på plats i dag är mer stabil och säker , tack vare våra framgångar med att bekämpa terrorismen " , sade han .
Regeringen fortsätter att bygga upp de områden som har förstörts av terrorister , för att återupprätta normaliteten .
Det finns nu alla förutsättningar för frivilligt återvändande av flyktingar till landet de tvingades lämna på grund av terrorism och unilaterala ekonomiska åtgärder som riktades mot deras dagliga liv och uppehälle .
FN uppskattar att mer än 5,5 miljoner syrier har flytt landet sedan kriget började 2011 .
Ytterligare sex miljoner människor som fortfarande bor i landet har behov av humanitärt stöd .
Enligt Al @-@ Moualem skulle den syriska regimen välkomna hjälp att återuppbygga det förstörda landet .
Men han betonade att den inte tar emot villkorat stöd eller hjälp från länder som har stöttat upproret .
Europa avgick med segern i Ryder Cup i Paris
Team Europa har vunnit 2018 års Ryder Cup genom att besegra Team USA med slutställningen 16,5 mot 10,5 vid Le Golf National utanför Paris i Frankrike .
USA har nu förlorat sex gånger i rad på europeisk mark och har inte vunnit Ryder Cup i Europa sedan 1993 .
Europa vann igen när den danske kaptenen Thomas Bjørns team uppnådde de 14,5 poäng som krävdes för att slå USA .
Den amerikanska stjärnan Phil Mickelson , som fick kämpa hårt under större delen av turneringen , hamnade i vattnet vid utslaget på det 16:e hålets par 3 @-@ bana , och förlorade mot Francesco Molinari .
Den italienske golfspelaren Molinari glänste i alla rundor och blev en av fyra spelare som någonsin har gjort 5 @-@ 0 @-@ 0 sedan turneringens nuvarande format infördes 1979 .
Amerikanen Jordan Spieth slogs ut 5 & 4 av det europeiska lagets lägst rankade spelare , Thorbjørn Olesen från Danmark .
Världens högst rankade spelare , Dustin Johnson , föll 2 & 1 mot Ian Poulter från England , som kan ha gjort sin sista Ryder Cup .
Spanjoren Sergio Garcia , som är en veteran med åtta Ryder Cup bakom sig , blev turneringens mest framgångsrika europé någonsin med 25,5 karriärpoäng .
" Jag brukar inte gråta , men i dag kan jag inte hjälpa det .
Det har varit ett tufft år .
Jag är så tacksam för att Thomas valde mig och trodde på mig .
Jag är så glad , så glad att vinna tillbaka segern .
Det handlar om laget , och jag är glad att jag kunde vara till hjälp " , sade en rörd Garcia efter Europalagets seger .
Han lämnade över stafettpinnen till sin landsman John Ram som besegrade den amerikanska golflegenden Tiger Woods 2 & 1 i singel på söndagen .
" Vilken otrolig stolthet , att få slå Tiger Woods . Jag är uppvuxen med att titta på honom , , sade den 23 @-@ årige Rahm .
Woods förlorade alla sina fyra matcher i Frankrike , och har nu resultatet 13 @-@ 21 @-@ 3 för sin karriär i Ryder cup .
En besynnerlig statistik för en av världens bästa spelare någonsin , som har vunnit 14 majortitlar , vilket endast har överträffats av Jack Nicklaus .
Team USA kämpade hela helgen med att hitta fairway , med undantag för Patrick Reed , Justin Thomas och Tony Finau , som spelade högklassig golf under hela turneringen .
Den amerikanske kaptenen Jim Furyk sade efter lagets nedslående prestation : " Jag är stolt över de här killarna , de har kämpat .
Det var dags i morse när vi höjde temperaturen i Europa .
Vi tog fajten .
Hatten av för Thomas .
Han är en fantastisk kapten .
Alla hans 12 spelare spelade riktigt bra .
Vi ska omgruppera oss , jag ska arbeta med USA:s PGA @-@ tour och vår Ryder Cup @-@ kommitté och så går vi vidare .
Jag älskar de här 12 killarna och är stolt över att vara kapten .
Man får buga och bocka .
De spelade bättre än vi " .
Algblomningen : Halterna minskar i Pinellas , Manatee och Sarasota
Den senaste rapporten från Floridas fiske- och viltkommission visar en generell minskning i koncentrationer av algblomning för delar av området runt Tampa Bay .
Enligt kommissionen rapporteras ojämnare blomningar i områdena runt storkommunerna Pinellas , Manatee , Sarasota , Charlotte och Collier . Detta kan tyda på minskade halter .
Algblomningen sträcker sig längs drygt 20 mil av kusten , från norra Pinellas till södra Lee .
Fläckar kan ses ungefär en och en halv mil ut i havet utanför storkommunen Hillsborough , men på färre platser jämfört med förra veckan .
Algblomning har också observerats i storkommunen Pasco .
Medelhöga koncentrationer i eller utanför kusten i Pinellas har rapporterats under den gångna veckan . Utanför Hillsboroughs kust låga till höga koncentrationer , bakgrundskoncentrationer till höga koncentrationer i Manatee , bakgrundskoncentrationer till höga koncentrationer i eller utanför kusten i Sarasota , bakgrundskoncentrationer till medelhöga koncentrationer i eller utanför kusten i Lee , och låga koncentrationer i Collier .
Rapporter om andningsirritation fortsätter att komma från storkommunerna Pinellas , Manatee , Sarasota , Lee och Collier .
Det förekom inga rapporter om andningsirritation i nordvästra Florida den gångna veckan .
