version https://git-lfs.github.com/spec/v1
oid sha256:f5d6946d22efaa4a31751aa9aa262cbfca12ad236331f5f76cb592fd0c2f902b
size 155590080
